//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.08.2021 21:35:32
// Design Name: 
// Module Name: Activation_Rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module Activation_Rom(
  input load_mem
);
    reg [31:0] mem [511:0];
    always @(posedge load_mem)
    begin
        mem[0] = 32'b00000000000001011100000000000001;
        mem[1] = 32'b00000000000001011100000000000001;
        mem[2] = 32'b00000000000001101100000000000001;
        mem[3] = 32'b00000000000001101100000000000001;
        mem[4] = 32'b00000000000001101100000000000001;
        mem[5] = 32'b00000000000001101100000000000001;
        mem[6] = 32'b00000000000001101100000000000001;
        mem[7] = 32'b00000000000001111100000000000001;
        mem[8] = 32'b00000000000001111100000000000001;
        mem[9] = 32'b00000000000001111100000000000001;
        mem[10] = 32'b00000000000001111100000000000001;
        mem[11] = 32'b00000000000001111100000000000001;
        mem[12] = 32'b00000000000010001100000000000001;
        mem[13] = 32'b00000000000010001100000000000001;
        mem[14] = 32'b00000000000010001100000000000001;
        mem[15] = 32'b00000000000010011100000000000001;
        mem[16] = 32'b00000000000010011100000000000001;
        mem[17] = 32'b00000000000010011100000000000001;
        mem[18] = 32'b00000000000010011100000000000001;
        mem[19] = 32'b00000000000010101100000000000001;
        mem[20] = 32'b00000000000010101100000000000001;
        mem[21] = 32'b00000000000010101100000000000001;
        mem[22] = 32'b00000000000010111100000000000001;
        mem[23] = 32'b00000000000010111100000000000001;
        mem[24] = 32'b00000000000010111100000000000001;
        mem[25] = 32'b00000000000011001100000000000001;
        mem[26] = 32'b00000000000011001100000000000001;
        mem[27] = 32'b00000000000011011100000000000001;
        mem[28] = 32'b00000000000011011100000000000001;
        mem[29] = 32'b00000000000011101100000000000001;
        mem[30] = 32'b00000000000011101100000000000001;
        mem[31] = 32'b00000000000011101100000000000001;
        mem[32] = 32'b00000000000011111100000000000001;
        mem[33] = 32'b00000000000011111100000000000001;
        mem[34] = 32'b00000000000100001100000000000001;
        mem[35] = 32'b00000000000100001100000000000001;
        mem[36] = 32'b00000000000100011100000000000001;
        mem[37] = 32'b00000000000100101100000000000001;
        mem[38] = 32'b00000000000100101100000000000001;
        mem[39] = 32'b00000000000100111100000000000001;
        mem[40] = 32'b00000000000100111100000000000001;
        mem[41] = 32'b00000000000101001100000000000001;
        mem[42] = 32'b00000000000101011100000000000001;
        mem[43] = 32'b00000000000101011100000000000001;
        mem[44] = 32'b00000000000101101100000000000001;
        mem[45] = 32'b00000000000101111100000000000001;
        mem[46] = 32'b00000000000101111100000000000001;
        mem[47] = 32'b00000000000110001100000000000001;
        mem[48] = 32'b00000000000110011100000000000001;
        mem[49] = 32'b00000000000110101100000000000001;
        mem[50] = 32'b00000000000110111100000000000001;
        mem[51] = 32'b00000000000110111100000000000001;
        mem[52] = 32'b00000000000111001100000000000001;
        mem[53] = 32'b00000000000111011100000000000001;
        mem[54] = 32'b00000000000111101100000000000001;
        mem[55] = 32'b00000000000111111100000000000001;
        mem[56] = 32'b00000000001000001100000000000001;
        mem[57] = 32'b00000000001000011100000000000001;
        mem[58] = 32'b00000000001000101100000000000001;
        mem[59] = 32'b00000000001000111100000000000001;
        mem[60] = 32'b00000000001001001100000000000001;
        mem[61] = 32'b00000000001001101100000000000001;
        mem[62] = 32'b00000000001001111100000000000001;
        mem[63] = 32'b00000000001010001100000000000001;
        mem[64] = 32'b00000000001010011100000000000001;
        mem[65] = 32'b00000000001010111100000000000001;
        mem[66] = 32'b00000000001011001100000000000001;
        mem[67] = 32'b00000000001011011100000000000001;
        mem[68] = 32'b00000000001011111100000000000001;
        mem[69] = 32'b00000000001100001100000000000001;
        mem[70] = 32'b00000000001100101100000000000001;
        mem[71] = 32'b00000000001100111100000000000001;
        mem[72] = 32'b00000000001101011100000000000001;
        mem[73] = 32'b00000000001101111100000000000001;
        mem[74] = 32'b00000000001110011100000000000001;
        mem[75] = 32'b00000000001110101100000000000001;
        mem[76] = 32'b00000000001111001100000000000001;
        mem[77] = 32'b00000000001111101100000000000001;
        mem[78] = 32'b00000000010000001100000000000001;
        mem[79] = 32'b00000000010000101100000000000001;
        mem[80] = 32'b00000000010001001100000000000001;
        mem[81] = 32'b00000000010001101100000000000001;
        mem[82] = 32'b00000000010010011100000000000001;
        mem[83] = 32'b00000000010010111100000000000001;
        mem[84] = 32'b00000000010011011100000000000001;
        mem[85] = 32'b00000000010100001100000000000001;
        mem[86] = 32'b00000000010100101100000000000001;
        mem[87] = 32'b00000000010101011100000000000001;
        mem[88] = 32'b00000000010110001100000000000001;
        mem[89] = 32'b00000000010110111100000000000010;
        mem[90] = 32'b00000000010111011100000000000010;
        mem[91] = 32'b00000000011000001100000000000010;
        mem[92] = 32'b00000000011000111100000000000010;
        mem[93] = 32'b00000000011001111100000000000010;
        mem[94] = 32'b00000000011010101100000000000010;
        mem[95] = 32'b00000000011011011100000000000010;
        mem[96] = 32'b00000000011100011100000000000010;
        mem[97] = 32'b00000000011101001100000000000010;
        mem[98] = 32'b00000000011110001100000000000010;
        mem[99] = 32'b00000000011111001100000000000010;
        mem[100] = 32'b00000000100000001100000000000011;
        mem[101] = 32'b00000000100001001100000000000011;
        mem[102] = 32'b00000000100010001100000000000011;
        mem[103] = 32'b00000000100011001100000000000011;
        mem[104] = 32'b00000000100100001100000000000011;
        mem[105] = 32'b00000000100101011100000000000011;
        mem[106] = 32'b00000000100110101100000000000011;
        mem[107] = 32'b00000000100111111100000000000100;
        mem[108] = 32'b00000000101001001100000000000100;
        mem[109] = 32'b00000000101010011100000000000100;
        mem[110] = 32'b00000000101011101100000000000100;
        mem[111] = 32'b00000000101101001100000000000101;
        mem[112] = 32'b00000000101110011100000000000101;
        mem[113] = 32'b00000000101111111100000000000101;
        mem[114] = 32'b00000000110001011100000000000101;
        mem[115] = 32'b00000000110010111100000000000110;
        mem[116] = 32'b00000000110100101100000000000110;
        mem[117] = 32'b00000000110110001100000000000110;
        mem[118] = 32'b00000000110111111100000000000111;
        mem[119] = 32'b00000000111001101100000000000111;
        mem[120] = 32'b00000000111011011100000000001000;
        mem[121] = 32'b00000000111101011100000000001000;
        mem[122] = 32'b00000000111111001100000000001001;
        mem[123] = 32'b00000001000001001100000000001001;
        mem[124] = 32'b00000001000011001100000000001010;
        mem[125] = 32'b00000001000101011100000000001010;
        mem[126] = 32'b00000001000111011100000000001011;
        mem[127] = 32'b00000001001001101100000000001011;
        mem[128] = 32'b00000001001011111100000000001100;
        mem[129] = 32'b00000001001110011100000000001101;
        mem[130] = 32'b00000001010000111100000000001110;
        mem[131] = 32'b00000001010011011100000000001111;
        mem[132] = 32'b00000001010101111100000000010000;
        mem[133] = 32'b00000001011000101100000000010000;
        mem[134] = 32'b00000001011011011100000000010010;
        mem[135] = 32'b00000001011110001100000000010011;
        mem[136] = 32'b00000001100001001100000000010100;
        mem[137] = 32'b00000001100100001100000000010101;
        mem[138] = 32'b00000001100111001100000000010110;
        mem[139] = 32'b00000001101010011100000000011000;
        mem[140] = 32'b00000001101101101100000000011001;
        mem[141] = 32'b00000001110000111100000000011011;
        mem[142] = 32'b00000001110100011100000000011101;
        mem[143] = 32'b00000001111000001100000000011110;
        mem[144] = 32'b00000001111011111100000000100000;
        mem[145] = 32'b00000001111111101100000000100010;
        mem[146] = 32'b00000010000011011100000000100101;
        mem[147] = 32'b00000010000111101100000000100111;
        mem[148] = 32'b00000010001011101100000000101001;
        mem[149] = 32'b00000010001111111100000000101100;
        mem[150] = 32'b00000010010100011100000000101111;
        mem[151] = 32'b00000010011000111100000000110010;
        mem[152] = 32'b00000010011101101100000000110101;
        mem[153] = 32'b00000010100010011100000000111000;
        mem[154] = 32'b00000010100111011100000000111100;
        mem[155] = 32'b00000010101100011100000001000000;
        mem[156] = 32'b00000010110001101100000001000100;
        mem[157] = 32'b00000010110111001100000001001000;
        mem[158] = 32'b00000010111100101100000001001101;
        mem[159] = 32'b00000011000010011100000001010010;
        mem[160] = 32'b00000011001000001100000001010111;
        mem[161] = 32'b00000011001110001100000001011100;
        mem[162] = 32'b00000011010100011100000001100010;
        mem[163] = 32'b00000011011010101100000001101000;
        mem[164] = 32'b00000011100001011100000001101111;
        mem[165] = 32'b00000011101000001100000001110110;
        mem[166] = 32'b00000011101110111100000001111110;
        mem[167] = 32'b00000011110110001100000010000110;
        mem[168] = 32'b00000011111101011100000010001110;
        mem[169] = 32'b00000100000100111100000010011000;
        mem[170] = 32'b00000100001100101100000010100001;
        mem[171] = 32'b00000100010100101100000010101100;
        mem[172] = 32'b00000100011100111100000010110111;
        mem[173] = 32'b00000100100101001100000011000010;
        mem[174] = 32'b00000100101101111100000011001111;
        mem[175] = 32'b00000100110110101100000011011100;
        mem[176] = 32'b00000100111111111100000011101010;
        mem[177] = 32'b00000101001001001100000011111001;
        mem[178] = 32'b00000101010010101100000100001001;
        mem[179] = 32'b00000101011100101100000100011010;
        mem[180] = 32'b00000101100110101100000100101100;
        mem[181] = 32'b00000101110001001100000100111111;
        mem[182] = 32'b00000101111011101100000101010011;
        mem[183] = 32'b00000110000110101100000101101001;
        mem[184] = 32'b00000110010001101100000101111111;
        mem[185] = 32'b00000110011101001100000110011000;
        mem[186] = 32'b00000110101000111100000110110010;
        mem[187] = 32'b00000110110101001100000111001101;
        mem[188] = 32'b00000111000001011100000111101011;
        mem[189] = 32'b00000111001110001100001000001010;
        mem[190] = 32'b00000111011010111100001000101011;
        mem[191] = 32'b00000111101000011100001001001110;
        mem[192] = 32'b00000111110101111100001001110011;
        mem[193] = 32'b00001000000011111100001010011011;
        mem[194] = 32'b00001000010010001100001011000101;
        mem[195] = 32'b00001000100000101100001011110001;
        mem[196] = 32'b00001000101111101100001100100001;
        mem[197] = 32'b00001000111110111100001101010011;
        mem[198] = 32'b00001001001110011100001110001000;
        mem[199] = 32'b00001001011110011100001111000001;
        mem[200] = 32'b00001001101110101100001111111101;
        mem[201] = 32'b00001001111111011100010000111101;
        mem[202] = 32'b00001010010000011100010010000000;
        mem[203] = 32'b00001010100001111100010011001000;
        mem[204] = 32'b00001010110011101100010100010011;
        mem[205] = 32'b00001011000101111100010101100100;
        mem[206] = 32'b00001011011000011100010110111001;
        mem[207] = 32'b00001011101011001100011000010011;
        mem[208] = 32'b00001011111110011100011001110010;
        mem[209] = 32'b00001100010010001100011011010110;
        mem[210] = 32'b00001100100110001100011101000001;
        mem[211] = 32'b00001100111010101100011110110001;
        mem[212] = 32'b00001101001111011100100000101000;
        mem[213] = 32'b00001101100100101100100010100110;
        mem[214] = 32'b00001101111010001100100100101010;
        mem[215] = 32'b00001110010000001100100110110110;
        mem[216] = 32'b00001110100110101100101001001010;
        mem[217] = 32'b00001110111101011100101011100101;
        mem[218] = 32'b00001111010100011100101110001001;
        mem[219] = 32'b00001111101011111100110000110101;
        mem[220] = 32'b00010000000011101100110011101010;
        mem[221] = 32'b00010000011011111100110110101001;
        mem[222] = 32'b00010000110100101100111001110001;
        mem[223] = 32'b00010001001101101100111101000011;
        mem[224] = 32'b00010001100110111101000000011111;
        mem[225] = 32'b00010010000000101101000100000101;
        mem[226] = 32'b00010010011010101101000111110111;
        mem[227] = 32'b00010010110101001101001011110100;
        mem[228] = 32'b00010011001111111101001111111100;
        mem[229] = 32'b00010011101010111101010100001111;
        mem[230] = 32'b00010100000110011101011000101111;
        mem[231] = 32'b00010100100010001101011101011010;
        mem[232] = 32'b00010100111110001101100010010010;
        mem[233] = 32'b00010101011010011101100111010110;
        mem[234] = 32'b00010101110111001101101100100110;
        mem[235] = 32'b00010110010100001101110010000010;
        mem[236] = 32'b00010110110001011101110111101011;
        mem[237] = 32'b00010111001110101101111101011111;
        mem[238] = 32'b00010111101100011110000011100000;
        mem[239] = 32'b00011000001010011110001001101101;
        mem[240] = 32'b00011000101000101110010000000110;
        mem[241] = 32'b00011001000111001110010110101001;
        mem[242] = 32'b00011001100101101110011101011000;
        mem[243] = 32'b00011010000100011110100100010001;
        mem[244] = 32'b00011010100011011110101011010100;
        mem[245] = 32'b00011011000010101110110010100001;
        mem[246] = 32'b00011011100001111110111001110110;
        mem[247] = 32'b00011100000001011111000001010100;
        mem[248] = 32'b00011100100000111111001000111001;
        mem[249] = 32'b00011101000000101111010000100100;
        mem[250] = 32'b00011101100000011111011000010101;
        mem[251] = 32'b00011110000000001111100000001011;
        mem[252] = 32'b00011110100000001111101000000101;
        mem[253] = 32'b00011111000000001111110000000010;
        mem[254] = 32'b00011111100000001111111000000001;
        mem[255] = 32'b00100000000000000000000000000000;
        mem[256] = 32'b00100000011111110000000111111111;
        mem[257] = 32'b00100000111111110000001111111110;
        mem[258] = 32'b00100001011111110000010111111011;
        mem[259] = 32'b00100001111111110000011111110101;
        mem[260] = 32'b00100010011111100000100111101011;
        mem[261] = 32'b00100010111111010000101111011100;
        mem[262] = 32'b00100011011111000000110111000111;
        mem[263] = 32'b00100011111110100000111110101100;
        mem[264] = 32'b00100100011110000001000110001010;
        mem[265] = 32'b00100100111101010001001101011111;
        mem[266] = 32'b00100101011100100001010100101100;
        mem[267] = 32'b00100101111011100001011011101111;
        mem[268] = 32'b00100110011010010001100010101000;
        mem[269] = 32'b00100110111000110001101001010111;
        mem[270] = 32'b00100111010111010001101111111010;
        mem[271] = 32'b00100111110101100001110110010011;
        mem[272] = 32'b00101000010011100001111100100000;
        mem[273] = 32'b00101000110001010010000010100001;
        mem[274] = 32'b00101001001110100010001000010101;
        mem[275] = 32'b00101001101011110010001101111110;
        mem[276] = 32'b00101010001000110010010011011010;
        mem[277] = 32'b00101010100101100010011000101010;
        mem[278] = 32'b00101011000001110010011101101110;
        mem[279] = 32'b00101011011101110010100010100110;
        mem[280] = 32'b00101011111001100010100111010001;
        mem[281] = 32'b00101100010101000010101011110001;
        mem[282] = 32'b00101100110000000010110000000100;
        mem[283] = 32'b00101101001010110010110100001100;
        mem[284] = 32'b00101101100101010010111000001001;
        mem[285] = 32'b00101101111111010010111011111011;
        mem[286] = 32'b00101110011001000010111111100001;
        mem[287] = 32'b00101110110010010011000010111101;
        mem[288] = 32'b00101111001011010011000110001111;
        mem[289] = 32'b00101111100100000011001001010111;
        mem[290] = 32'b00101111111100010011001100010110;
        mem[291] = 32'b00110000010100000011001111001011;
        mem[292] = 32'b00110000101011100011010001110111;
        mem[293] = 32'b00110001000010100011010100011011;
        mem[294] = 32'b00110001011001010011010110110110;
        mem[295] = 32'b00110001101111110011011001001010;
        mem[296] = 32'b00110010000101110011011011010110;
        mem[297] = 32'b00110010011011010011011101011010;
        mem[298] = 32'b00110010110000100011011111011000;
        mem[299] = 32'b00110011000101010011100001001111;
        mem[300] = 32'b00110011011001110011100010111111;
        mem[301] = 32'b00110011101101110011100100101010;
        mem[302] = 32'b00110100000001100011100110001110;
        mem[303] = 32'b00110100010100110011100111101101;
        mem[304] = 32'b00110100100111100011101001000111;
        mem[305] = 32'b00110100111010000011101010011100;
        mem[306] = 32'b00110101001100010011101011101101;
        mem[307] = 32'b00110101011110000011101100111000;
        mem[308] = 32'b00110101101111100011101110000000;
        mem[309] = 32'b00110110000000100011101111000011;
        mem[310] = 32'b00110110010001010011110000000011;
        mem[311] = 32'b00110110100001100011110000111111;
        mem[312] = 32'b00110110110001100011110001111000;
        mem[313] = 32'b00110111000001000011110010101101;
        mem[314] = 32'b00110111010000010011110011011111;
        mem[315] = 32'b00110111011111010011110100001111;
        mem[316] = 32'b00110111101101110011110100111011;
        mem[317] = 32'b00110111111100000011110101100101;
        mem[318] = 32'b00111000001010000011110110001101;
        mem[319] = 32'b00111000010111100011110110110010;
        mem[320] = 32'b00111000100101000011110111010101;
        mem[321] = 32'b00111000110001110011110111110110;
        mem[322] = 32'b00111000111110100011111000010101;
        mem[323] = 32'b00111001001010110011111000110011;
        mem[324] = 32'b00111001010111000011111001001110;
        mem[325] = 32'b00111001100010110011111001101000;
        mem[326] = 32'b00111001101110010011111010000001;
        mem[327] = 32'b00111001111001010011111010010111;
        mem[328] = 32'b00111010000100010011111010101101;
        mem[329] = 32'b00111010001110110011111011000001;
        mem[330] = 32'b00111010011001010011111011010100;
        mem[331] = 32'b00111010100011010011111011100110;
        mem[332] = 32'b00111010101101010011111011110111;
        mem[333] = 32'b00111010110110110011111100000111;
        mem[334] = 32'b00111011000000000011111100010110;
        mem[335] = 32'b00111011001001010011111100100100;
        mem[336] = 32'b00111011010010000011111100110001;
        mem[337] = 32'b00111011011010110011111100111110;
        mem[338] = 32'b00111011100011000011111101001001;
        mem[339] = 32'b00111011101011010011111101010100;
        mem[340] = 32'b00111011110011010011111101011111;
        mem[341] = 32'b00111011111011000011111101101000;
        mem[342] = 32'b00111100000010100011111101110010;
        mem[343] = 32'b00111100001001110011111101111010;
        mem[344] = 32'b00111100010001000011111110000010;
        mem[345] = 32'b00111100010111110011111110001010;
        mem[346] = 32'b00111100011110100011111110010001;
        mem[347] = 32'b00111100100101010011111110011000;
        mem[348] = 32'b00111100101011100011111110011110;
        mem[349] = 32'b00111100110001110011111110100100;
        mem[350] = 32'b00111100110111110011111110101001;
        mem[351] = 32'b00111100111101100011111110101110;
        mem[352] = 32'b00111101000011010011111110110011;
        mem[353] = 32'b00111101001000110011111110111000;
        mem[354] = 32'b00111101001110010011111110111100;
        mem[355] = 32'b00111101010011100011111111000000;
        mem[356] = 32'b00111101011000100011111111000100;
        mem[357] = 32'b00111101011101100011111111001000;
        mem[358] = 32'b00111101100010010011111111001011;
        mem[359] = 32'b00111101100111000011111111001110;
        mem[360] = 32'b00111101101011100011111111010001;
        mem[361] = 32'b00111101110000000011111111010100;
        mem[362] = 32'b00111101110100010011111111010111;
        mem[363] = 32'b00111101111000010011111111011001;
        mem[364] = 32'b00111101111100100011111111011011;
        mem[365] = 32'b00111110000000010011111111011110;
        mem[366] = 32'b00111110000100000011111111100000;
        mem[367] = 32'b00111110000111110011111111100010;
        mem[368] = 32'b00111110001011100011111111100011;
        mem[369] = 32'b00111110001111000011111111100101;
        mem[370] = 32'b00111110010010010011111111100111;
        mem[371] = 32'b00111110010101100011111111101000;
        mem[372] = 32'b00111110011000110011111111101010;
        mem[373] = 32'b00111110011011110011111111101011;
        mem[374] = 32'b00111110011110110011111111101100;
        mem[375] = 32'b00111110100001110011111111101101;
        mem[376] = 32'b00111110100100100011111111101110;
        mem[377] = 32'b00111110100111010011111111110000;
        mem[378] = 32'b00111110101010000011111111110000;
        mem[379] = 32'b00111110101100100011111111110001;
        mem[380] = 32'b00111110101111000011111111110010;
        mem[381] = 32'b00111110110001100011111111110011;
        mem[382] = 32'b00111110110100000011111111110100;
        mem[383] = 32'b00111110110110010011111111110101;
        mem[384] = 32'b00111110111000100011111111110101;
        mem[385] = 32'b00111110111010100011111111110110;
        mem[386] = 32'b00111110111100110011111111110110;
        mem[387] = 32'b00111110111110110011111111110111;
        mem[388] = 32'b00111111000000110011111111110111;
        mem[389] = 32'b00111111000010100011111111111000;
        mem[390] = 32'b00111111000100100011111111111000;
        mem[391] = 32'b00111111000110010011111111111001;
        mem[392] = 32'b00111111001000000011111111111001;
        mem[393] = 32'b00111111001001110011111111111010;
        mem[394] = 32'b00111111001011010011111111111010;
        mem[395] = 32'b00111111001101000011111111111010;
        mem[396] = 32'b00111111001110100011111111111011;
        mem[397] = 32'b00111111010000000011111111111011;
        mem[398] = 32'b00111111010001100011111111111011;
        mem[399] = 32'b00111111010010110011111111111011;
        mem[400] = 32'b00111111010100010011111111111100;
        mem[401] = 32'b00111111010101100011111111111100;
        mem[402] = 32'b00111111010110110011111111111100;
        mem[403] = 32'b00111111011000000011111111111100;
        mem[404] = 32'b00111111011001010011111111111101;
        mem[405] = 32'b00111111011010100011111111111101;
        mem[406] = 32'b00111111011011110011111111111101;
        mem[407] = 32'b00111111011100110011111111111101;
        mem[408] = 32'b00111111011101110011111111111101;
        mem[409] = 32'b00111111011110110011111111111101;
        mem[410] = 32'b00111111011111110011111111111101;
        mem[411] = 32'b00111111100000110011111111111110;
        mem[412] = 32'b00111111100001110011111111111110;
        mem[413] = 32'b00111111100010110011111111111110;
        mem[414] = 32'b00111111100011100011111111111110;
        mem[415] = 32'b00111111100100100011111111111110;
        mem[416] = 32'b00111111100101010011111111111110;
        mem[417] = 32'b00111111100110000011111111111110;
        mem[418] = 32'b00111111100111000011111111111110;
        mem[419] = 32'b00111111100111110011111111111110;
        mem[420] = 32'b00111111101000100011111111111110;
        mem[421] = 32'b00111111101001000011111111111110;
        mem[422] = 32'b00111111101001110011111111111111;
        mem[423] = 32'b00111111101010100011111111111111;
        mem[424] = 32'b00111111101011010011111111111111;
        mem[425] = 32'b00111111101011110011111111111111;
        mem[426] = 32'b00111111101100100011111111111111;
        mem[427] = 32'b00111111101101000011111111111111;
        mem[428] = 32'b00111111101101100011111111111111;
        mem[429] = 32'b00111111101110010011111111111111;
        mem[430] = 32'b00111111101110110011111111111111;
        mem[431] = 32'b00111111101111010011111111111111;
        mem[432] = 32'b00111111101111110011111111111111;
        mem[433] = 32'b00111111110000010011111111111111;
        mem[434] = 32'b00111111110000110011111111111111;
        mem[435] = 32'b00111111110001010011111111111111;
        mem[436] = 32'b00111111110001100011111111111111;
        mem[437] = 32'b00111111110010000011111111111111;
        mem[438] = 32'b00111111110010100011111111111111;
        mem[439] = 32'b00111111110011000011111111111111;
        mem[440] = 32'b00111111110011010011111111111111;
        mem[441] = 32'b00111111110011110011111111111111;
        mem[442] = 32'b00111111110100000011111111111111;
        mem[443] = 32'b00111111110100100011111111111111;
        mem[444] = 32'b00111111110100110011111111111111;
        mem[445] = 32'b00111111110101000011111111111111;
        mem[446] = 32'b00111111110101100011111111111111;
        mem[447] = 32'b00111111110101110011111111111111;
        mem[448] = 32'b00111111110110000011111111111111;
        mem[449] = 32'b00111111110110010011111111111111;
        mem[450] = 32'b00111111110110110011111111111111;
        mem[451] = 32'b00111111110111000011111111111111;
        mem[452] = 32'b00111111110111010011111111111111;
        mem[453] = 32'b00111111110111100011111111111111;
        mem[454] = 32'b00111111110111110011111111111111;
        mem[455] = 32'b00111111111000000011111111111111;
        mem[456] = 32'b00111111111000010011111111111111;
        mem[457] = 32'b00111111111000100011111111111111;
        mem[458] = 32'b00111111111000110011111111111111;
        mem[459] = 32'b00111111111001000011111111111111;
        mem[460] = 32'b00111111111001000011111111111111;
        mem[461] = 32'b00111111111001010011111111111111;
        mem[462] = 32'b00111111111001100011111111111111;
        mem[463] = 32'b00111111111001110011111111111111;
        mem[464] = 32'b00111111111010000011111111111111;
        mem[465] = 32'b00111111111010000011111111111111;
        mem[466] = 32'b00111111111010010011111111111111;
        mem[467] = 32'b00111111111010100011111111111111;
        mem[468] = 32'b00111111111010100011111111111111;
        mem[469] = 32'b00111111111010110011111111111111;
        mem[470] = 32'b00111111111011000011111111111111;
        mem[471] = 32'b00111111111011000011111111111111;
        mem[472] = 32'b00111111111011010011111111111111;
        mem[473] = 32'b00111111111011010011111111111111;
        mem[474] = 32'b00111111111011100011111111111111;
        mem[475] = 32'b00111111111011110011111111111111;
        mem[476] = 32'b00111111111011110011111111111111;
        mem[477] = 32'b00111111111100000011111111111111;
        mem[478] = 32'b00111111111100000011111111111111;
        mem[479] = 32'b00111111111100010011111111111111;
        mem[480] = 32'b00111111111100010011111111111111;
        mem[481] = 32'b00111111111100010011111111111111;
        mem[482] = 32'b00111111111100100011111111111111;
        mem[483] = 32'b00111111111100100011111111111111;
        mem[484] = 32'b00111111111100110011111111111111;
        mem[485] = 32'b00111111111100110011111111111111;
        mem[486] = 32'b00111111111101000011111111111111;
        mem[487] = 32'b00111111111101000011111111111111;
        mem[488] = 32'b00111111111101000011111111111111;
        mem[489] = 32'b00111111111101010011111111111111;
        mem[490] = 32'b00111111111101010011111111111111;
        mem[491] = 32'b00111111111101010011111111111111;
        mem[492] = 32'b00111111111101100011111111111111;
        mem[493] = 32'b00111111111101100011111111111111;
        mem[494] = 32'b00111111111101100011111111111111;
        mem[495] = 32'b00111111111101100011111111111111;
        mem[496] = 32'b00111111111101110011111111111111;
        mem[497] = 32'b00111111111101110011111111111111;
        mem[498] = 32'b00111111111101110011111111111111;
        mem[499] = 32'b00111111111110000011111111111111;
        mem[500] = 32'b00111111111110000011111111111111;
        mem[501] = 32'b00111111111110000011111111111111;
        mem[502] = 32'b00111111111110000011111111111111;
        mem[503] = 32'b00111111111110000011111111111111;
        mem[504] = 32'b00111111111110010011111111111111;
        mem[505] = 32'b00111111111110010011111111111111;
        mem[506] = 32'b00111111111110010011111111111111;
        mem[507] = 32'b00111111111110010011111111111111;
        mem[508] = 32'b00111111111110010011111111111111;
        mem[509] = 32'b00111111111110100011111111111111;
        mem[510] = 32'b00111111111110100011111111111111;
    end
endmodule