//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.08.2021 21:35:32
// Design Name: 
// Module Name: Activation_Rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Activation_Rom(
  input load_mem
);
    reg [31:0] mem [1023:0];
    always @(posedge load_mem)
    begin
        mem[0] = 32'b00000000000000001100000000000001;
        mem[1] = 32'b00000000000000001100000000000001;
        mem[2] = 32'b00000000000000001100000000000001;
        mem[3] = 32'b00000000000000001100000000000001;
        mem[4] = 32'b00000000000000001100000000000001;
        mem[5] = 32'b00000000000000001100000000000001;
        mem[6] = 32'b00000000000000001100000000000001;
        mem[7] = 32'b00000000000000001100000000000001;
        mem[8] = 32'b00000000000000001100000000000001;
        mem[9] = 32'b00000000000000001100000000000001;
        mem[10] = 32'b00000000000000001100000000000001;
        mem[11] = 32'b00000000000000001100000000000001;
        mem[12] = 32'b00000000000000001100000000000001;
        mem[13] = 32'b00000000000000001100000000000001;
        mem[14] = 32'b00000000000000001100000000000001;
        mem[15] = 32'b00000000000000001100000000000001;
        mem[16] = 32'b00000000000000001100000000000001;
        mem[17] = 32'b00000000000000001100000000000001;
        mem[18] = 32'b00000000000000001100000000000001;
        mem[19] = 32'b00000000000000001100000000000001;
        mem[20] = 32'b00000000000000001100000000000001;
        mem[21] = 32'b00000000000000001100000000000001;
        mem[22] = 32'b00000000000000001100000000000001;
        mem[23] = 32'b00000000000000001100000000000001;
        mem[24] = 32'b00000000000000001100000000000001;
        mem[25] = 32'b00000000000000001100000000000001;
        mem[26] = 32'b00000000000000001100000000000001;
        mem[27] = 32'b00000000000000001100000000000001;
        mem[28] = 32'b00000000000000001100000000000001;
        mem[29] = 32'b00000000000000001100000000000001;
        mem[30] = 32'b00000000000000001100000000000001;
        mem[31] = 32'b00000000000000001100000000000001;
        mem[32] = 32'b00000000000000001100000000000001;
        mem[33] = 32'b00000000000000001100000000000001;
        mem[34] = 32'b00000000000000001100000000000001;
        mem[35] = 32'b00000000000000001100000000000001;
        mem[36] = 32'b00000000000000001100000000000001;
        mem[37] = 32'b00000000000000001100000000000001;
        mem[38] = 32'b00000000000000001100000000000001;
        mem[39] = 32'b00000000000000001100000000000001;
        mem[40] = 32'b00000000000000001100000000000001;
        mem[41] = 32'b00000000000000001100000000000001;
        mem[42] = 32'b00000000000000001100000000000001;
        mem[43] = 32'b00000000000000001100000000000001;
        mem[44] = 32'b00000000000000001100000000000001;
        mem[45] = 32'b00000000000000001100000000000001;
        mem[46] = 32'b00000000000000001100000000000001;
        mem[47] = 32'b00000000000000001100000000000001;
        mem[48] = 32'b00000000000000001100000000000001;
        mem[49] = 32'b00000000000000001100000000000001;
        mem[50] = 32'b00000000000000001100000000000001;
        mem[51] = 32'b00000000000000001100000000000001;
        mem[52] = 32'b00000000000000001100000000000001;
        mem[53] = 32'b00000000000000001100000000000001;
        mem[54] = 32'b00000000000000001100000000000001;
        mem[55] = 32'b00000000000000001100000000000001;
        mem[56] = 32'b00000000000000001100000000000001;
        mem[57] = 32'b00000000000000001100000000000001;
        mem[58] = 32'b00000000000000001100000000000001;
        mem[59] = 32'b00000000000000001100000000000001;
        mem[60] = 32'b00000000000000001100000000000001;
        mem[61] = 32'b00000000000000001100000000000001;
        mem[62] = 32'b00000000000000001100000000000001;
        mem[63] = 32'b00000000000000001100000000000001;
        mem[64] = 32'b00000000000000001100000000000001;
        mem[65] = 32'b00000000000000001100000000000001;
        mem[66] = 32'b00000000000000001100000000000001;
        mem[67] = 32'b00000000000000001100000000000001;
        mem[68] = 32'b00000000000000001100000000000001;
        mem[69] = 32'b00000000000000001100000000000001;
        mem[70] = 32'b00000000000000001100000000000001;
        mem[71] = 32'b00000000000000001100000000000001;
        mem[72] = 32'b00000000000000001100000000000001;
        mem[73] = 32'b00000000000000001100000000000001;
        mem[74] = 32'b00000000000000001100000000000001;
        mem[75] = 32'b00000000000000001100000000000001;
        mem[76] = 32'b00000000000000001100000000000001;
        mem[77] = 32'b00000000000000001100000000000001;
        mem[78] = 32'b00000000000000001100000000000001;
        mem[79] = 32'b00000000000000001100000000000001;
        mem[80] = 32'b00000000000000001100000000000001;
        mem[81] = 32'b00000000000000001100000000000001;
        mem[82] = 32'b00000000000000001100000000000001;
        mem[83] = 32'b00000000000000001100000000000001;
        mem[84] = 32'b00000000000000001100000000000001;
        mem[85] = 32'b00000000000000001100000000000001;
        mem[86] = 32'b00000000000000001100000000000001;
        mem[87] = 32'b00000000000000001100000000000001;
        mem[88] = 32'b00000000000000001100000000000001;
        mem[89] = 32'b00000000000000001100000000000001;
        mem[90] = 32'b00000000000000001100000000000001;
        mem[91] = 32'b00000000000000001100000000000001;
        mem[92] = 32'b00000000000000001100000000000001;
        mem[93] = 32'b00000000000000001100000000000001;
        mem[94] = 32'b00000000000000001100000000000001;
        mem[95] = 32'b00000000000000001100000000000001;
        mem[96] = 32'b00000000000000001100000000000001;
        mem[97] = 32'b00000000000000001100000000000001;
        mem[98] = 32'b00000000000000001100000000000001;
        mem[99] = 32'b00000000000000001100000000000001;
        mem[100] = 32'b00000000000000001100000000000001;
        mem[101] = 32'b00000000000000001100000000000001;
        mem[102] = 32'b00000000000000001100000000000001;
        mem[103] = 32'b00000000000000001100000000000001;
        mem[104] = 32'b00000000000000001100000000000001;
        mem[105] = 32'b00000000000000001100000000000001;
        mem[106] = 32'b00000000000000001100000000000001;
        mem[107] = 32'b00000000000000001100000000000001;
        mem[108] = 32'b00000000000000001100000000000001;
        mem[109] = 32'b00000000000000001100000000000001;
        mem[110] = 32'b00000000000000001100000000000001;
        mem[111] = 32'b00000000000000001100000000000001;
        mem[112] = 32'b00000000000000001100000000000001;
        mem[113] = 32'b00000000000000001100000000000001;
        mem[114] = 32'b00000000000000001100000000000001;
        mem[115] = 32'b00000000000000001100000000000001;
        mem[116] = 32'b00000000000000001100000000000001;
        mem[117] = 32'b00000000000000001100000000000001;
        mem[118] = 32'b00000000000000001100000000000001;
        mem[119] = 32'b00000000000000001100000000000001;
        mem[120] = 32'b00000000000000001100000000000001;
        mem[121] = 32'b00000000000000001100000000000001;
        mem[122] = 32'b00000000000000001100000000000001;
        mem[123] = 32'b00000000000000001100000000000001;
        mem[124] = 32'b00000000000000001100000000000001;
        mem[125] = 32'b00000000000000001100000000000001;
        mem[126] = 32'b00000000000000001100000000000001;
        mem[127] = 32'b00000000000000001100000000000001;
        mem[128] = 32'b00000000000000001100000000000001;
        mem[129] = 32'b00000000000000001100000000000001;
        mem[130] = 32'b00000000000000001100000000000001;
        mem[131] = 32'b00000000000000001100000000000001;
        mem[132] = 32'b00000000000000001100000000000001;
        mem[133] = 32'b00000000000000001100000000000001;
        mem[134] = 32'b00000000000000001100000000000001;
        mem[135] = 32'b00000000000000001100000000000001;
        mem[136] = 32'b00000000000000001100000000000001;
        mem[137] = 32'b00000000000000001100000000000001;
        mem[138] = 32'b00000000000000001100000000000001;
        mem[139] = 32'b00000000000000001100000000000001;
        mem[140] = 32'b00000000000000001100000000000001;
        mem[141] = 32'b00000000000000001100000000000001;
        mem[142] = 32'b00000000000000001100000000000001;
        mem[143] = 32'b00000000000000001100000000000001;
        mem[144] = 32'b00000000000000001100000000000001;
        mem[145] = 32'b00000000000000001100000000000001;
        mem[146] = 32'b00000000000000001100000000000001;
        mem[147] = 32'b00000000000000001100000000000001;
        mem[148] = 32'b00000000000000001100000000000001;
        mem[149] = 32'b00000000000000001100000000000001;
        mem[150] = 32'b00000000000000001100000000000001;
        mem[151] = 32'b00000000000000001100000000000001;
        mem[152] = 32'b00000000000000001100000000000001;
        mem[153] = 32'b00000000000000001100000000000001;
        mem[154] = 32'b00000000000000001100000000000001;
        mem[155] = 32'b00000000000000001100000000000001;
        mem[156] = 32'b00000000000000001100000000000001;
        mem[157] = 32'b00000000000000001100000000000001;
        mem[158] = 32'b00000000000000001100000000000001;
        mem[159] = 32'b00000000000000001100000000000001;
        mem[160] = 32'b00000000000000001100000000000001;
        mem[161] = 32'b00000000000000001100000000000001;
        mem[162] = 32'b00000000000000001100000000000001;
        mem[163] = 32'b00000000000000001100000000000001;
        mem[164] = 32'b00000000000000001100000000000001;
        mem[165] = 32'b00000000000000001100000000000001;
        mem[166] = 32'b00000000000000001100000000000001;
        mem[167] = 32'b00000000000000001100000000000001;
        mem[168] = 32'b00000000000000001100000000000001;
        mem[169] = 32'b00000000000000001100000000000001;
        mem[170] = 32'b00000000000000001100000000000001;
        mem[171] = 32'b00000000000000001100000000000001;
        mem[172] = 32'b00000000000000001100000000000001;
        mem[173] = 32'b00000000000000001100000000000001;
        mem[174] = 32'b00000000000000001100000000000001;
        mem[175] = 32'b00000000000000001100000000000001;
        mem[176] = 32'b00000000000000001100000000000001;
        mem[177] = 32'b00000000000000001100000000000001;
        mem[178] = 32'b00000000000000001100000000000001;
        mem[179] = 32'b00000000000000001100000000000001;
        mem[180] = 32'b00000000000000001100000000000001;
        mem[181] = 32'b00000000000000001100000000000001;
        mem[182] = 32'b00000000000000001100000000000001;
        mem[183] = 32'b00000000000000001100000000000001;
        mem[184] = 32'b00000000000000001100000000000001;
        mem[185] = 32'b00000000000000001100000000000001;
        mem[186] = 32'b00000000000000001100000000000001;
        mem[187] = 32'b00000000000000001100000000000001;
        mem[188] = 32'b00000000000000001100000000000001;
        mem[189] = 32'b00000000000000001100000000000001;
        mem[190] = 32'b00000000000000001100000000000001;
        mem[191] = 32'b00000000000000001100000000000001;
        mem[192] = 32'b00000000000000001100000000000001;
        mem[193] = 32'b00000000000000001100000000000001;
        mem[194] = 32'b00000000000000001100000000000001;
        mem[195] = 32'b00000000000000001100000000000001;
        mem[196] = 32'b00000000000000001100000000000001;
        mem[197] = 32'b00000000000000001100000000000001;
        mem[198] = 32'b00000000000000001100000000000001;
        mem[199] = 32'b00000000000000001100000000000001;
        mem[200] = 32'b00000000000000001100000000000001;
        mem[201] = 32'b00000000000000011100000000000001;
        mem[202] = 32'b00000000000000011100000000000001;
        mem[203] = 32'b00000000000000011100000000000001;
        mem[204] = 32'b00000000000000011100000000000001;
        mem[205] = 32'b00000000000000011100000000000001;
        mem[206] = 32'b00000000000000011100000000000001;
        mem[207] = 32'b00000000000000011100000000000001;
        mem[208] = 32'b00000000000000011100000000000001;
        mem[209] = 32'b00000000000000011100000000000001;
        mem[210] = 32'b00000000000000011100000000000001;
        mem[211] = 32'b00000000000000011100000000000001;
        mem[212] = 32'b00000000000000011100000000000001;
        mem[213] = 32'b00000000000000011100000000000001;
        mem[214] = 32'b00000000000000011100000000000001;
        mem[215] = 32'b00000000000000011100000000000001;
        mem[216] = 32'b00000000000000011100000000000001;
        mem[217] = 32'b00000000000000011100000000000001;
        mem[218] = 32'b00000000000000011100000000000001;
        mem[219] = 32'b00000000000000011100000000000001;
        mem[220] = 32'b00000000000000011100000000000001;
        mem[221] = 32'b00000000000000011100000000000001;
        mem[222] = 32'b00000000000000011100000000000001;
        mem[223] = 32'b00000000000000101100000000000001;
        mem[224] = 32'b00000000000000101100000000000001;
        mem[225] = 32'b00000000000000101100000000000001;
        mem[226] = 32'b00000000000000101100000000000001;
        mem[227] = 32'b00000000000000101100000000000001;
        mem[228] = 32'b00000000000000101100000000000001;
        mem[229] = 32'b00000000000000101100000000000001;
        mem[230] = 32'b00000000000000101100000000000001;
        mem[231] = 32'b00000000000000101100000000000001;
        mem[232] = 32'b00000000000000101100000000000001;
        mem[233] = 32'b00000000000000101100000000000001;
        mem[234] = 32'b00000000000000101100000000000001;
        mem[235] = 32'b00000000000000101100000000000001;
        mem[236] = 32'b00000000000000111100000000000001;
        mem[237] = 32'b00000000000000111100000000000001;
        mem[238] = 32'b00000000000000111100000000000001;
        mem[239] = 32'b00000000000000111100000000000001;
        mem[240] = 32'b00000000000000111100000000000001;
        mem[241] = 32'b00000000000000111100000000000001;
        mem[242] = 32'b00000000000000111100000000000001;
        mem[243] = 32'b00000000000000111100000000000001;
        mem[244] = 32'b00000000000000111100000000000001;
        mem[245] = 32'b00000000000001001100000000000001;
        mem[246] = 32'b00000000000001001100000000000001;
        mem[247] = 32'b00000000000001001100000000000001;
        mem[248] = 32'b00000000000001001100000000000001;
        mem[249] = 32'b00000000000001001100000000000001;
        mem[250] = 32'b00000000000001001100000000000001;
        mem[251] = 32'b00000000000001001100000000000001;
        mem[252] = 32'b00000000000001011100000000000001;
        mem[253] = 32'b00000000000001011100000000000001;
        mem[254] = 32'b00000000000001011100000000000001;
        mem[255] = 32'b00000000000001011100000000000001;
        mem[256] = 32'b00000000000001011100000000000001;
        mem[257] = 32'b00000000000001011100000000000001;
        mem[258] = 32'b00000000000001101100000000000001;
        mem[259] = 32'b00000000000001101100000000000001;
        mem[260] = 32'b00000000000001101100000000000001;
        mem[261] = 32'b00000000000001101100000000000001;
        mem[262] = 32'b00000000000001101100000000000001;
        mem[263] = 32'b00000000000001111100000000000001;
        mem[264] = 32'b00000000000001111100000000000001;
        mem[265] = 32'b00000000000001111100000000000001;
        mem[266] = 32'b00000000000001111100000000000001;
        mem[267] = 32'b00000000000001111100000000000001;
        mem[268] = 32'b00000000000010001100000000000001;
        mem[269] = 32'b00000000000010001100000000000001;
        mem[270] = 32'b00000000000010001100000000000001;
        mem[271] = 32'b00000000000010011100000000000001;
        mem[272] = 32'b00000000000010011100000000000001;
        mem[273] = 32'b00000000000010011100000000000001;
        mem[274] = 32'b00000000000010011100000000000001;
        mem[275] = 32'b00000000000010101100000000000001;
        mem[276] = 32'b00000000000010101100000000000001;
        mem[277] = 32'b00000000000010101100000000000001;
        mem[278] = 32'b00000000000010111100000000000001;
        mem[279] = 32'b00000000000010111100000000000001;
        mem[280] = 32'b00000000000010111100000000000001;
        mem[281] = 32'b00000000000011001100000000000001;
        mem[282] = 32'b00000000000011001100000000000001;
        mem[283] = 32'b00000000000011011100000000000001;
        mem[284] = 32'b00000000000011011100000000000001;
        mem[285] = 32'b00000000000011101100000000000001;
        mem[286] = 32'b00000000000011101100000000000001;
        mem[287] = 32'b00000000000011101100000000000001;
        mem[288] = 32'b00000000000011111100000000000001;
        mem[289] = 32'b00000000000011111100000000000001;
        mem[290] = 32'b00000000000100001100000000000001;
        mem[291] = 32'b00000000000100001100000000000001;
        mem[292] = 32'b00000000000100011100000000000001;
        mem[293] = 32'b00000000000100101100000000000001;
        mem[294] = 32'b00000000000100101100000000000001;
        mem[295] = 32'b00000000000100111100000000000001;
        mem[296] = 32'b00000000000100111100000000000001;
        mem[297] = 32'b00000000000101001100000000000001;
        mem[298] = 32'b00000000000101011100000000000001;
        mem[299] = 32'b00000000000101011100000000000001;
        mem[300] = 32'b00000000000101101100000000000001;
        mem[301] = 32'b00000000000101111100000000000001;
        mem[302] = 32'b00000000000101111100000000000001;
        mem[303] = 32'b00000000000110001100000000000001;
        mem[304] = 32'b00000000000110011100000000000001;
        mem[305] = 32'b00000000000110101100000000000001;
        mem[306] = 32'b00000000000110111100000000000001;
        mem[307] = 32'b00000000000110111100000000000001;
        mem[308] = 32'b00000000000111001100000000000001;
        mem[309] = 32'b00000000000111011100000000000001;
        mem[310] = 32'b00000000000111101100000000000001;
        mem[311] = 32'b00000000000111111100000000000001;
        mem[312] = 32'b00000000001000001100000000000001;
        mem[313] = 32'b00000000001000011100000000000001;
        mem[314] = 32'b00000000001000101100000000000001;
        mem[315] = 32'b00000000001000111100000000000001;
        mem[316] = 32'b00000000001001001100000000000001;
        mem[317] = 32'b00000000001001101100000000000001;
        mem[318] = 32'b00000000001001111100000000000001;
        mem[319] = 32'b00000000001010001100000000000001;
        mem[320] = 32'b00000000001010011100000000000001;
        mem[321] = 32'b00000000001010111100000000000001;
        mem[322] = 32'b00000000001011001100000000000001;
        mem[323] = 32'b00000000001011011100000000000001;
        mem[324] = 32'b00000000001011111100000000000001;
        mem[325] = 32'b00000000001100001100000000000001;
        mem[326] = 32'b00000000001100101100000000000001;
        mem[327] = 32'b00000000001100111100000000000001;
        mem[328] = 32'b00000000001101011100000000000001;
        mem[329] = 32'b00000000001101111100000000000001;
        mem[330] = 32'b00000000001110011100000000000001;
        mem[331] = 32'b00000000001110101100000000000001;
        mem[332] = 32'b00000000001111001100000000000001;
        mem[333] = 32'b00000000001111101100000000000001;
        mem[334] = 32'b00000000010000001100000000000001;
        mem[335] = 32'b00000000010000101100000000000001;
        mem[336] = 32'b00000000010001001100000000000001;
        mem[337] = 32'b00000000010001101100000000000001;
        mem[338] = 32'b00000000010010011100000000000001;
        mem[339] = 32'b00000000010010111100000000000001;
        mem[340] = 32'b00000000010011011100000000000001;
        mem[341] = 32'b00000000010100001100000000000001;
        mem[342] = 32'b00000000010100101100000000000001;
        mem[343] = 32'b00000000010101011100000000000001;
        mem[344] = 32'b00000000010110001100000000000001;
        mem[345] = 32'b00000000010110111100000000000010;
        mem[346] = 32'b00000000010111011100000000000010;
        mem[347] = 32'b00000000011000001100000000000010;
        mem[348] = 32'b00000000011000111100000000000010;
        mem[349] = 32'b00000000011001111100000000000010;
        mem[350] = 32'b00000000011010101100000000000010;
        mem[351] = 32'b00000000011011011100000000000010;
        mem[352] = 32'b00000000011100011100000000000010;
        mem[353] = 32'b00000000011101001100000000000010;
        mem[354] = 32'b00000000011110001100000000000010;
        mem[355] = 32'b00000000011111001100000000000010;
        mem[356] = 32'b00000000100000001100000000000011;
        mem[357] = 32'b00000000100001001100000000000011;
        mem[358] = 32'b00000000100010001100000000000011;
        mem[359] = 32'b00000000100011001100000000000011;
        mem[360] = 32'b00000000100100001100000000000011;
        mem[361] = 32'b00000000100101011100000000000011;
        mem[362] = 32'b00000000100110101100000000000011;
        mem[363] = 32'b00000000100111111100000000000100;
        mem[364] = 32'b00000000101001001100000000000100;
        mem[365] = 32'b00000000101010011100000000000100;
        mem[366] = 32'b00000000101011101100000000000100;
        mem[367] = 32'b00000000101101001100000000000101;
        mem[368] = 32'b00000000101110011100000000000101;
        mem[369] = 32'b00000000101111111100000000000101;
        mem[370] = 32'b00000000110001011100000000000101;
        mem[371] = 32'b00000000110010111100000000000110;
        mem[372] = 32'b00000000110100101100000000000110;
        mem[373] = 32'b00000000110110001100000000000110;
        mem[374] = 32'b00000000110111111100000000000111;
        mem[375] = 32'b00000000111001101100000000000111;
        mem[376] = 32'b00000000111011011100000000001000;
        mem[377] = 32'b00000000111101011100000000001000;
        mem[378] = 32'b00000000111111001100000000001001;
        mem[379] = 32'b00000001000001001100000000001001;
        mem[380] = 32'b00000001000011001100000000001010;
        mem[381] = 32'b00000001000101011100000000001010;
        mem[382] = 32'b00000001000111011100000000001011;
        mem[383] = 32'b00000001001001101100000000001011;
        mem[384] = 32'b00000001001011111100000000001100;
        mem[385] = 32'b00000001001110011100000000001101;
        mem[386] = 32'b00000001010000111100000000001110;
        mem[387] = 32'b00000001010011011100000000001111;
        mem[388] = 32'b00000001010101111100000000010000;
        mem[389] = 32'b00000001011000101100000000010000;
        mem[390] = 32'b00000001011011011100000000010010;
        mem[391] = 32'b00000001011110001100000000010011;
        mem[392] = 32'b00000001100001001100000000010100;
        mem[393] = 32'b00000001100100001100000000010101;
        mem[394] = 32'b00000001100111001100000000010110;
        mem[395] = 32'b00000001101010011100000000011000;
        mem[396] = 32'b00000001101101101100000000011001;
        mem[397] = 32'b00000001110000111100000000011011;
        mem[398] = 32'b00000001110100011100000000011101;
        mem[399] = 32'b00000001111000001100000000011110;
        mem[400] = 32'b00000001111011111100000000100000;
        mem[401] = 32'b00000001111111101100000000100010;
        mem[402] = 32'b00000010000011011100000000100101;
        mem[403] = 32'b00000010000111101100000000100111;
        mem[404] = 32'b00000010001011101100000000101001;
        mem[405] = 32'b00000010001111111100000000101100;
        mem[406] = 32'b00000010010100011100000000101111;
        mem[407] = 32'b00000010011000111100000000110010;
        mem[408] = 32'b00000010011101101100000000110101;
        mem[409] = 32'b00000010100010011100000000111000;
        mem[410] = 32'b00000010100111011100000000111100;
        mem[411] = 32'b00000010101100011100000001000000;
        mem[412] = 32'b00000010110001101100000001000100;
        mem[413] = 32'b00000010110111001100000001001000;
        mem[414] = 32'b00000010111100101100000001001101;
        mem[415] = 32'b00000011000010011100000001010010;
        mem[416] = 32'b00000011001000001100000001010111;
        mem[417] = 32'b00000011001110001100000001011100;
        mem[418] = 32'b00000011010100011100000001100010;
        mem[419] = 32'b00000011011010101100000001101000;
        mem[420] = 32'b00000011100001011100000001101111;
        mem[421] = 32'b00000011101000001100000001110110;
        mem[422] = 32'b00000011101110111100000001111110;
        mem[423] = 32'b00000011110110001100000010000110;
        mem[424] = 32'b00000011111101011100000010001110;
        mem[425] = 32'b00000100000100111100000010011000;
        mem[426] = 32'b00000100001100101100000010100001;
        mem[427] = 32'b00000100010100101100000010101100;
        mem[428] = 32'b00000100011100111100000010110111;
        mem[429] = 32'b00000100100101001100000011000010;
        mem[430] = 32'b00000100101101111100000011001111;
        mem[431] = 32'b00000100110110101100000011011100;
        mem[432] = 32'b00000100111111111100000011101010;
        mem[433] = 32'b00000101001001001100000011111001;
        mem[434] = 32'b00000101010010101100000100001001;
        mem[435] = 32'b00000101011100101100000100011010;
        mem[436] = 32'b00000101100110101100000100101100;
        mem[437] = 32'b00000101110001001100000100111111;
        mem[438] = 32'b00000101111011101100000101010011;
        mem[439] = 32'b00000110000110101100000101101001;
        mem[440] = 32'b00000110010001101100000101111111;
        mem[441] = 32'b00000110011101001100000110011000;
        mem[442] = 32'b00000110101000111100000110110010;
        mem[443] = 32'b00000110110101001100000111001101;
        mem[444] = 32'b00000111000001011100000111101011;
        mem[445] = 32'b00000111001110001100001000001010;
        mem[446] = 32'b00000111011010111100001000101011;
        mem[447] = 32'b00000111101000011100001001001110;
        mem[448] = 32'b00000111110101111100001001110011;
        mem[449] = 32'b00001000000011111100001010011011;
        mem[450] = 32'b00001000010010001100001011000101;
        mem[451] = 32'b00001000100000101100001011110001;
        mem[452] = 32'b00001000101111101100001100100001;
        mem[453] = 32'b00001000111110111100001101010011;
        mem[454] = 32'b00001001001110011100001110001000;
        mem[455] = 32'b00001001011110011100001111000001;
        mem[456] = 32'b00001001101110101100001111111101;
        mem[457] = 32'b00001001111111011100010000111101;
        mem[458] = 32'b00001010010000011100010010000000;
        mem[459] = 32'b00001010100001111100010011001000;
        mem[460] = 32'b00001010110011101100010100010011;
        mem[461] = 32'b00001011000101111100010101100100;
        mem[462] = 32'b00001011011000011100010110111001;
        mem[463] = 32'b00001011101011001100011000010011;
        mem[464] = 32'b00001011111110011100011001110010;
        mem[465] = 32'b00001100010010001100011011010110;
        mem[466] = 32'b00001100100110001100011101000001;
        mem[467] = 32'b00001100111010101100011110110001;
        mem[468] = 32'b00001101001111011100100000101000;
        mem[469] = 32'b00001101100100101100100010100110;
        mem[470] = 32'b00001101111010001100100100101010;
        mem[471] = 32'b00001110010000001100100110110110;
        mem[472] = 32'b00001110100110101100101001001010;
        mem[473] = 32'b00001110111101011100101011100101;
        mem[474] = 32'b00001111010100011100101110001001;
        mem[475] = 32'b00001111101011111100110000110101;
        mem[476] = 32'b00010000000011101100110011101010;
        mem[477] = 32'b00010000011011111100110110101001;
        mem[478] = 32'b00010000110100101100111001110001;
        mem[479] = 32'b00010001001101101100111101000011;
        mem[480] = 32'b00010001100110111101000000011111;
        mem[481] = 32'b00010010000000101101000100000101;
        mem[482] = 32'b00010010011010101101000111110111;
        mem[483] = 32'b00010010110101001101001011110100;
        mem[484] = 32'b00010011001111111101001111111100;
        mem[485] = 32'b00010011101010111101010100001111;
        mem[486] = 32'b00010100000110011101011000101111;
        mem[487] = 32'b00010100100010001101011101011010;
        mem[488] = 32'b00010100111110001101100010010010;
        mem[489] = 32'b00010101011010011101100111010110;
        mem[490] = 32'b00010101110111001101101100100110;
        mem[491] = 32'b00010110010100001101110010000010;
        mem[492] = 32'b00010110110001011101110111101011;
        mem[493] = 32'b00010111001110101101111101011111;
        mem[494] = 32'b00010111101100011110000011100000;
        mem[495] = 32'b00011000001010011110001001101101;
        mem[496] = 32'b00011000101000101110010000000110;
        mem[497] = 32'b00011001000111001110010110101001;
        mem[498] = 32'b00011001100101101110011101011000;
        mem[499] = 32'b00011010000100011110100100010001;
        mem[500] = 32'b00011010100011011110101011010100;
        mem[501] = 32'b00011011000010101110110010100001;
        mem[502] = 32'b00011011100001111110111001110110;
        mem[503] = 32'b00011100000001011111000001010100;
        mem[504] = 32'b00011100100000111111001000111001;
        mem[505] = 32'b00011101000000101111010000100100;
        mem[506] = 32'b00011101100000011111011000010101;
        mem[507] = 32'b00011110000000001111100000001011;
        mem[508] = 32'b00011110100000001111101000000101;
        mem[509] = 32'b00011111000000001111110000000010;
        mem[510] = 32'b00011111100000001111111000000001;
        mem[511] = 32'b00100000000000000000000000000000;
        mem[512] = 32'b00100000011111110000000111111111;
        mem[513] = 32'b00100000111111110000001111111110;
        mem[514] = 32'b00100001011111110000010111111011;
        mem[515] = 32'b00100001111111110000011111110101;
        mem[516] = 32'b00100010011111100000100111101011;
        mem[517] = 32'b00100010111111010000101111011100;
        mem[518] = 32'b00100011011111000000110111000111;
        mem[519] = 32'b00100011111110100000111110101100;
        mem[520] = 32'b00100100011110000001000110001010;
        mem[521] = 32'b00100100111101010001001101011111;
        mem[522] = 32'b00100101011100100001010100101100;
        mem[523] = 32'b00100101111011100001011011101111;
        mem[524] = 32'b00100110011010010001100010101000;
        mem[525] = 32'b00100110111000110001101001010111;
        mem[526] = 32'b00100111010111010001101111111010;
        mem[527] = 32'b00100111110101100001110110010011;
        mem[528] = 32'b00101000010011100001111100100000;
        mem[529] = 32'b00101000110001010010000010100001;
        mem[530] = 32'b00101001001110100010001000010101;
        mem[531] = 32'b00101001101011110010001101111110;
        mem[532] = 32'b00101010001000110010010011011010;
        mem[533] = 32'b00101010100101100010011000101010;
        mem[534] = 32'b00101011000001110010011101101110;
        mem[535] = 32'b00101011011101110010100010100110;
        mem[536] = 32'b00101011111001100010100111010001;
        mem[537] = 32'b00101100010101000010101011110001;
        mem[538] = 32'b00101100110000000010110000000100;
        mem[539] = 32'b00101101001010110010110100001100;
        mem[540] = 32'b00101101100101010010111000001001;
        mem[541] = 32'b00101101111111010010111011111011;
        mem[542] = 32'b00101110011001000010111111100001;
        mem[543] = 32'b00101110110010010011000010111101;
        mem[544] = 32'b00101111001011010011000110001111;
        mem[545] = 32'b00101111100100000011001001010111;
        mem[546] = 32'b00101111111100010011001100010110;
        mem[547] = 32'b00110000010100000011001111001011;
        mem[548] = 32'b00110000101011100011010001110111;
        mem[549] = 32'b00110001000010100011010100011011;
        mem[550] = 32'b00110001011001010011010110110110;
        mem[551] = 32'b00110001101111110011011001001010;
        mem[552] = 32'b00110010000101110011011011010110;
        mem[553] = 32'b00110010011011010011011101011010;
        mem[554] = 32'b00110010110000100011011111011000;
        mem[555] = 32'b00110011000101010011100001001111;
        mem[556] = 32'b00110011011001110011100010111111;
        mem[557] = 32'b00110011101101110011100100101010;
        mem[558] = 32'b00110100000001100011100110001110;
        mem[559] = 32'b00110100010100110011100111101101;
        mem[560] = 32'b00110100100111100011101001000111;
        mem[561] = 32'b00110100111010000011101010011100;
        mem[562] = 32'b00110101001100010011101011101101;
        mem[563] = 32'b00110101011110000011101100111000;
        mem[564] = 32'b00110101101111100011101110000000;
        mem[565] = 32'b00110110000000100011101111000011;
        mem[566] = 32'b00110110010001010011110000000011;
        mem[567] = 32'b00110110100001100011110000111111;
        mem[568] = 32'b00110110110001100011110001111000;
        mem[569] = 32'b00110111000001000011110010101101;
        mem[570] = 32'b00110111010000010011110011011111;
        mem[571] = 32'b00110111011111010011110100001111;
        mem[572] = 32'b00110111101101110011110100111011;
        mem[573] = 32'b00110111111100000011110101100101;
        mem[574] = 32'b00111000001010000011110110001101;
        mem[575] = 32'b00111000010111100011110110110010;
        mem[576] = 32'b00111000100101000011110111010101;
        mem[577] = 32'b00111000110001110011110111110110;
        mem[578] = 32'b00111000111110100011111000010101;
        mem[579] = 32'b00111001001010110011111000110011;
        mem[580] = 32'b00111001010111000011111001001110;
        mem[581] = 32'b00111001100010110011111001101000;
        mem[582] = 32'b00111001101110010011111010000001;
        mem[583] = 32'b00111001111001010011111010010111;
        mem[584] = 32'b00111010000100010011111010101101;
        mem[585] = 32'b00111010001110110011111011000001;
        mem[586] = 32'b00111010011001010011111011010100;
        mem[587] = 32'b00111010100011010011111011100110;
        mem[588] = 32'b00111010101101010011111011110111;
        mem[589] = 32'b00111010110110110011111100000111;
        mem[590] = 32'b00111011000000000011111100010110;
        mem[591] = 32'b00111011001001010011111100100100;
        mem[592] = 32'b00111011010010000011111100110001;
        mem[593] = 32'b00111011011010110011111100111110;
        mem[594] = 32'b00111011100011000011111101001001;
        mem[595] = 32'b00111011101011010011111101010100;
        mem[596] = 32'b00111011110011010011111101011111;
        mem[597] = 32'b00111011111011000011111101101000;
        mem[598] = 32'b00111100000010100011111101110010;
        mem[599] = 32'b00111100001001110011111101111010;
        mem[600] = 32'b00111100010001000011111110000010;
        mem[601] = 32'b00111100010111110011111110001010;
        mem[602] = 32'b00111100011110100011111110010001;
        mem[603] = 32'b00111100100101010011111110011000;
        mem[604] = 32'b00111100101011100011111110011110;
        mem[605] = 32'b00111100110001110011111110100100;
        mem[606] = 32'b00111100110111110011111110101001;
        mem[607] = 32'b00111100111101100011111110101110;
        mem[608] = 32'b00111101000011010011111110110011;
        mem[609] = 32'b00111101001000110011111110111000;
        mem[610] = 32'b00111101001110010011111110111100;
        mem[611] = 32'b00111101010011100011111111000000;
        mem[612] = 32'b00111101011000100011111111000100;
        mem[613] = 32'b00111101011101100011111111001000;
        mem[614] = 32'b00111101100010010011111111001011;
        mem[615] = 32'b00111101100111000011111111001110;
        mem[616] = 32'b00111101101011100011111111010001;
        mem[617] = 32'b00111101110000000011111111010100;
        mem[618] = 32'b00111101110100010011111111010111;
        mem[619] = 32'b00111101111000010011111111011001;
        mem[620] = 32'b00111101111100100011111111011011;
        mem[621] = 32'b00111110000000010011111111011110;
        mem[622] = 32'b00111110000100000011111111100000;
        mem[623] = 32'b00111110000111110011111111100010;
        mem[624] = 32'b00111110001011100011111111100011;
        mem[625] = 32'b00111110001111000011111111100101;
        mem[626] = 32'b00111110010010010011111111100111;
        mem[627] = 32'b00111110010101100011111111101000;
        mem[628] = 32'b00111110011000110011111111101010;
        mem[629] = 32'b00111110011011110011111111101011;
        mem[630] = 32'b00111110011110110011111111101100;
        mem[631] = 32'b00111110100001110011111111101101;
        mem[632] = 32'b00111110100100100011111111101110;
        mem[633] = 32'b00111110100111010011111111110000;
        mem[634] = 32'b00111110101010000011111111110000;
        mem[635] = 32'b00111110101100100011111111110001;
        mem[636] = 32'b00111110101111000011111111110010;
        mem[637] = 32'b00111110110001100011111111110011;
        mem[638] = 32'b00111110110100000011111111110100;
        mem[639] = 32'b00111110110110010011111111110101;
        mem[640] = 32'b00111110111000100011111111110101;
        mem[641] = 32'b00111110111010100011111111110110;
        mem[642] = 32'b00111110111100110011111111110110;
        mem[643] = 32'b00111110111110110011111111110111;
        mem[644] = 32'b00111111000000110011111111110111;
        mem[645] = 32'b00111111000010100011111111111000;
        mem[646] = 32'b00111111000100100011111111111000;
        mem[647] = 32'b00111111000110010011111111111001;
        mem[648] = 32'b00111111001000000011111111111001;
        mem[649] = 32'b00111111001001110011111111111010;
        mem[650] = 32'b00111111001011010011111111111010;
        mem[651] = 32'b00111111001101000011111111111010;
        mem[652] = 32'b00111111001110100011111111111011;
        mem[653] = 32'b00111111010000000011111111111011;
        mem[654] = 32'b00111111010001100011111111111011;
        mem[655] = 32'b00111111010010110011111111111011;
        mem[656] = 32'b00111111010100010011111111111100;
        mem[657] = 32'b00111111010101100011111111111100;
        mem[658] = 32'b00111111010110110011111111111100;
        mem[659] = 32'b00111111011000000011111111111100;
        mem[660] = 32'b00111111011001010011111111111101;
        mem[661] = 32'b00111111011010100011111111111101;
        mem[662] = 32'b00111111011011110011111111111101;
        mem[663] = 32'b00111111011100110011111111111101;
        mem[664] = 32'b00111111011101110011111111111101;
        mem[665] = 32'b00111111011110110011111111111101;
        mem[666] = 32'b00111111011111110011111111111101;
        mem[667] = 32'b00111111100000110011111111111110;
        mem[668] = 32'b00111111100001110011111111111110;
        mem[669] = 32'b00111111100010110011111111111110;
        mem[670] = 32'b00111111100011100011111111111110;
        mem[671] = 32'b00111111100100100011111111111110;
        mem[672] = 32'b00111111100101010011111111111110;
        mem[673] = 32'b00111111100110000011111111111110;
        mem[674] = 32'b00111111100111000011111111111110;
        mem[675] = 32'b00111111100111110011111111111110;
        mem[676] = 32'b00111111101000100011111111111110;
        mem[677] = 32'b00111111101001000011111111111110;
        mem[678] = 32'b00111111101001110011111111111111;
        mem[679] = 32'b00111111101010100011111111111111;
        mem[680] = 32'b00111111101011010011111111111111;
        mem[681] = 32'b00111111101011110011111111111111;
        mem[682] = 32'b00111111101100100011111111111111;
        mem[683] = 32'b00111111101101000011111111111111;
        mem[684] = 32'b00111111101101100011111111111111;
        mem[685] = 32'b00111111101110010011111111111111;
        mem[686] = 32'b00111111101110110011111111111111;
        mem[687] = 32'b00111111101111010011111111111111;
        mem[688] = 32'b00111111101111110011111111111111;
        mem[689] = 32'b00111111110000010011111111111111;
        mem[690] = 32'b00111111110000110011111111111111;
        mem[691] = 32'b00111111110001010011111111111111;
        mem[692] = 32'b00111111110001100011111111111111;
        mem[693] = 32'b00111111110010000011111111111111;
        mem[694] = 32'b00111111110010100011111111111111;
        mem[695] = 32'b00111111110011000011111111111111;
        mem[696] = 32'b00111111110011010011111111111111;
        mem[697] = 32'b00111111110011110011111111111111;
        mem[698] = 32'b00111111110100000011111111111111;
        mem[699] = 32'b00111111110100100011111111111111;
        mem[700] = 32'b00111111110100110011111111111111;
        mem[701] = 32'b00111111110101000011111111111111;
        mem[702] = 32'b00111111110101100011111111111111;
        mem[703] = 32'b00111111110101110011111111111111;
        mem[704] = 32'b00111111110110000011111111111111;
        mem[705] = 32'b00111111110110010011111111111111;
        mem[706] = 32'b00111111110110110011111111111111;
        mem[707] = 32'b00111111110111000011111111111111;
        mem[708] = 32'b00111111110111010011111111111111;
        mem[709] = 32'b00111111110111100011111111111111;
        mem[710] = 32'b00111111110111110011111111111111;
        mem[711] = 32'b00111111111000000011111111111111;
        mem[712] = 32'b00111111111000010011111111111111;
        mem[713] = 32'b00111111111000100011111111111111;
        mem[714] = 32'b00111111111000110011111111111111;
        mem[715] = 32'b00111111111001000011111111111111;
        mem[716] = 32'b00111111111001000011111111111111;
        mem[717] = 32'b00111111111001010011111111111111;
        mem[718] = 32'b00111111111001100011111111111111;
        mem[719] = 32'b00111111111001110011111111111111;
        mem[720] = 32'b00111111111010000011111111111111;
        mem[721] = 32'b00111111111010000011111111111111;
        mem[722] = 32'b00111111111010010011111111111111;
        mem[723] = 32'b00111111111010100011111111111111;
        mem[724] = 32'b00111111111010100011111111111111;
        mem[725] = 32'b00111111111010110011111111111111;
        mem[726] = 32'b00111111111011000011111111111111;
        mem[727] = 32'b00111111111011000011111111111111;
        mem[728] = 32'b00111111111011010011111111111111;
        mem[729] = 32'b00111111111011010011111111111111;
        mem[730] = 32'b00111111111011100011111111111111;
        mem[731] = 32'b00111111111011110011111111111111;
        mem[732] = 32'b00111111111011110011111111111111;
        mem[733] = 32'b00111111111100000011111111111111;
        mem[734] = 32'b00111111111100000011111111111111;
        mem[735] = 32'b00111111111100010011111111111111;
        mem[736] = 32'b00111111111100010011111111111111;
        mem[737] = 32'b00111111111100010011111111111111;
        mem[738] = 32'b00111111111100100011111111111111;
        mem[739] = 32'b00111111111100100011111111111111;
        mem[740] = 32'b00111111111100110011111111111111;
        mem[741] = 32'b00111111111100110011111111111111;
        mem[742] = 32'b00111111111101000011111111111111;
        mem[743] = 32'b00111111111101000011111111111111;
        mem[744] = 32'b00111111111101000011111111111111;
        mem[745] = 32'b00111111111101010011111111111111;
        mem[746] = 32'b00111111111101010011111111111111;
        mem[747] = 32'b00111111111101010011111111111111;
        mem[748] = 32'b00111111111101100011111111111111;
        mem[749] = 32'b00111111111101100011111111111111;
        mem[750] = 32'b00111111111101100011111111111111;
        mem[751] = 32'b00111111111101100011111111111111;
        mem[752] = 32'b00111111111101110011111111111111;
        mem[753] = 32'b00111111111101110011111111111111;
        mem[754] = 32'b00111111111101110011111111111111;
        mem[755] = 32'b00111111111110000011111111111111;
        mem[756] = 32'b00111111111110000011111111111111;
        mem[757] = 32'b00111111111110000011111111111111;
        mem[758] = 32'b00111111111110000011111111111111;
        mem[759] = 32'b00111111111110000011111111111111;
        mem[760] = 32'b00111111111110010011111111111111;
        mem[761] = 32'b00111111111110010011111111111111;
        mem[762] = 32'b00111111111110010011111111111111;
        mem[763] = 32'b00111111111110010011111111111111;
        mem[764] = 32'b00111111111110010011111111111111;
        mem[765] = 32'b00111111111110100011111111111111;
        mem[766] = 32'b00111111111110100011111111111111;
        mem[767] = 32'b00111111111110100011111111111111;
        mem[768] = 32'b00111111111110100011111111111111;
        mem[769] = 32'b00111111111110100011111111111111;
        mem[770] = 32'b00111111111110100011111111111111;
        mem[771] = 32'b00111111111110110011111111111111;
        mem[772] = 32'b00111111111110110011111111111111;
        mem[773] = 32'b00111111111110110011111111111111;
        mem[774] = 32'b00111111111110110011111111111111;
        mem[775] = 32'b00111111111110110011111111111111;
        mem[776] = 32'b00111111111110110011111111111111;
        mem[777] = 32'b00111111111110110011111111111111;
        mem[778] = 32'b00111111111111000011111111111111;
        mem[779] = 32'b00111111111111000011111111111111;
        mem[780] = 32'b00111111111111000011111111111111;
        mem[781] = 32'b00111111111111000011111111111111;
        mem[782] = 32'b00111111111111000011111111111111;
        mem[783] = 32'b00111111111111000011111111111111;
        mem[784] = 32'b00111111111111000011111111111111;
        mem[785] = 32'b00111111111111000011111111111111;
        mem[786] = 32'b00111111111111000011111111111111;
        mem[787] = 32'b00111111111111010011111111111111;
        mem[788] = 32'b00111111111111010011111111111111;
        mem[789] = 32'b00111111111111010011111111111111;
        mem[790] = 32'b00111111111111010011111111111111;
        mem[791] = 32'b00111111111111010011111111111111;
        mem[792] = 32'b00111111111111010011111111111111;
        mem[793] = 32'b00111111111111010011111111111111;
        mem[794] = 32'b00111111111111010011111111111111;
        mem[795] = 32'b00111111111111010011111111111111;
        mem[796] = 32'b00111111111111010011111111111111;
        mem[797] = 32'b00111111111111010011111111111111;
        mem[798] = 32'b00111111111111010011111111111111;
        mem[799] = 32'b00111111111111010011111111111111;
        mem[800] = 32'b00111111111111100011111111111111;
        mem[801] = 32'b00111111111111100011111111111111;
        mem[802] = 32'b00111111111111100011111111111111;
        mem[803] = 32'b00111111111111100011111111111111;
        mem[804] = 32'b00111111111111100011111111111111;
        mem[805] = 32'b00111111111111100011111111111111;
        mem[806] = 32'b00111111111111100011111111111111;
        mem[807] = 32'b00111111111111100011111111111111;
        mem[808] = 32'b00111111111111100011111111111111;
        mem[809] = 32'b00111111111111100011111111111111;
        mem[810] = 32'b00111111111111100011111111111111;
        mem[811] = 32'b00111111111111100011111111111111;
        mem[812] = 32'b00111111111111100011111111111111;
        mem[813] = 32'b00111111111111100011111111111111;
        mem[814] = 32'b00111111111111100011111111111111;
        mem[815] = 32'b00111111111111100011111111111111;
        mem[816] = 32'b00111111111111100011111111111111;
        mem[817] = 32'b00111111111111100011111111111111;
        mem[818] = 32'b00111111111111100011111111111111;
        mem[819] = 32'b00111111111111100011111111111111;
        mem[820] = 32'b00111111111111100011111111111111;
        mem[821] = 32'b00111111111111100011111111111111;
        mem[822] = 32'b00111111111111110011111111111111;
        mem[823] = 32'b00111111111111110011111111111111;
        mem[824] = 32'b00111111111111110011111111111111;
        mem[825] = 32'b00111111111111110011111111111111;
        mem[826] = 32'b00111111111111110011111111111111;
        mem[827] = 32'b00111111111111110011111111111111;
        mem[828] = 32'b00111111111111110011111111111111;
        mem[829] = 32'b00111111111111110011111111111111;
        mem[830] = 32'b00111111111111110011111111111111;
        mem[831] = 32'b00111111111111110011111111111111;
        mem[832] = 32'b00111111111111110011111111111111;
        mem[833] = 32'b00111111111111110011111111111111;
        mem[834] = 32'b00111111111111110011111111111111;
        mem[835] = 32'b00111111111111110011111111111111;
        mem[836] = 32'b00111111111111110011111111111111;
        mem[837] = 32'b00111111111111110011111111111111;
        mem[838] = 32'b00111111111111110011111111111111;
        mem[839] = 32'b00111111111111110011111111111111;
        mem[840] = 32'b00111111111111110011111111111111;
        mem[841] = 32'b00111111111111110011111111111111;
        mem[842] = 32'b00111111111111110011111111111111;
        mem[843] = 32'b00111111111111110011111111111111;
        mem[844] = 32'b00111111111111110011111111111111;
        mem[845] = 32'b00111111111111110011111111111111;
        mem[846] = 32'b00111111111111110011111111111111;
        mem[847] = 32'b00111111111111110011111111111111;
        mem[848] = 32'b00111111111111110011111111111111;
        mem[849] = 32'b00111111111111110011111111111111;
        mem[850] = 32'b00111111111111110011111111111111;
        mem[851] = 32'b00111111111111110011111111111111;
        mem[852] = 32'b00111111111111110011111111111111;
        mem[853] = 32'b00111111111111110011111111111111;
        mem[854] = 32'b00111111111111110011111111111111;
        mem[855] = 32'b00111111111111110011111111111111;
        mem[856] = 32'b00111111111111110011111111111111;
        mem[857] = 32'b00111111111111110011111111111111;
        mem[858] = 32'b00111111111111110011111111111111;
        mem[859] = 32'b00111111111111110011111111111111;
        mem[860] = 32'b00111111111111110011111111111111;
        mem[861] = 32'b00111111111111110011111111111111;
        mem[862] = 32'b00111111111111110011111111111111;
        mem[863] = 32'b00111111111111110011111111111111;
        mem[864] = 32'b00111111111111110011111111111111;
        mem[865] = 32'b00111111111111110011111111111111;
        mem[866] = 32'b00111111111111110011111111111111;
        mem[867] = 32'b00111111111111110011111111111111;
        mem[868] = 32'b00111111111111110011111111111111;
        mem[869] = 32'b00111111111111110011111111111111;
        mem[870] = 32'b00111111111111110011111111111111;
        mem[871] = 32'b00111111111111110011111111111111;
        mem[872] = 32'b00111111111111110011111111111111;
        mem[873] = 32'b00111111111111110011111111111111;
        mem[874] = 32'b00111111111111110011111111111111;
        mem[875] = 32'b00111111111111110011111111111111;
        mem[876] = 32'b00111111111111110011111111111111;
        mem[877] = 32'b00111111111111110011111111111111;
        mem[878] = 32'b00111111111111110011111111111111;
        mem[879] = 32'b00111111111111110011111111111111;
        mem[880] = 32'b00111111111111110011111111111111;
        mem[881] = 32'b00111111111111110011111111111111;
        mem[882] = 32'b00111111111111110011111111111111;
        mem[883] = 32'b00111111111111110011111111111111;
        mem[884] = 32'b00111111111111110011111111111111;
        mem[885] = 32'b00111111111111110011111111111111;
        mem[886] = 32'b00111111111111110011111111111111;
        mem[887] = 32'b00111111111111110011111111111111;
        mem[888] = 32'b00111111111111110011111111111111;
        mem[889] = 32'b00111111111111110011111111111111;
        mem[890] = 32'b00111111111111110011111111111111;
        mem[891] = 32'b00111111111111110011111111111111;
        mem[892] = 32'b00111111111111110011111111111111;
        mem[893] = 32'b00111111111111110011111111111111;
        mem[894] = 32'b00111111111111110011111111111111;
        mem[895] = 32'b00111111111111110011111111111111;
        mem[896] = 32'b00111111111111110011111111111111;
        mem[897] = 32'b00111111111111110011111111111111;
        mem[898] = 32'b00111111111111110011111111111111;
        mem[899] = 32'b00111111111111110011111111111111;
        mem[900] = 32'b00111111111111110011111111111111;
        mem[901] = 32'b00111111111111110011111111111111;
        mem[902] = 32'b00111111111111110011111111111111;
        mem[903] = 32'b00111111111111110011111111111111;
        mem[904] = 32'b00111111111111110011111111111111;
        mem[905] = 32'b00111111111111110011111111111111;
        mem[906] = 32'b00111111111111110011111111111111;
        mem[907] = 32'b00111111111111110011111111111111;
        mem[908] = 32'b00111111111111110011111111111111;
        mem[909] = 32'b00111111111111110011111111111111;
        mem[910] = 32'b00111111111111110011111111111111;
        mem[911] = 32'b00111111111111110011111111111111;
        mem[912] = 32'b00111111111111110011111111111111;
        mem[913] = 32'b00111111111111110011111111111111;
        mem[914] = 32'b00111111111111110011111111111111;
        mem[915] = 32'b00111111111111110011111111111111;
        mem[916] = 32'b00111111111111110011111111111111;
        mem[917] = 32'b00111111111111110011111111111111;
        mem[918] = 32'b00111111111111110011111111111111;
        mem[919] = 32'b00111111111111110011111111111111;
        mem[920] = 32'b00111111111111110011111111111111;
        mem[921] = 32'b00111111111111110011111111111111;
        mem[922] = 32'b00111111111111110011111111111111;
        mem[923] = 32'b00111111111111110011111111111111;
        mem[924] = 32'b00111111111111110011111111111111;
        mem[925] = 32'b00111111111111110011111111111111;
        mem[926] = 32'b00111111111111110011111111111111;
        mem[927] = 32'b00111111111111110011111111111111;
        mem[928] = 32'b00111111111111110011111111111111;
        mem[929] = 32'b00111111111111110011111111111111;
        mem[930] = 32'b00111111111111110011111111111111;
        mem[931] = 32'b00111111111111110011111111111111;
        mem[932] = 32'b00111111111111110011111111111111;
        mem[933] = 32'b00111111111111110011111111111111;
        mem[934] = 32'b00111111111111110011111111111111;
        mem[935] = 32'b00111111111111110011111111111111;
        mem[936] = 32'b00111111111111110011111111111111;
        mem[937] = 32'b00111111111111110011111111111111;
        mem[938] = 32'b00111111111111110011111111111111;
        mem[939] = 32'b00111111111111110011111111111111;
        mem[940] = 32'b00111111111111110011111111111111;
        mem[941] = 32'b00111111111111110011111111111111;
        mem[942] = 32'b00111111111111110011111111111111;
        mem[943] = 32'b00111111111111110011111111111111;
        mem[944] = 32'b00111111111111110011111111111111;
        mem[945] = 32'b00111111111111110011111111111111;
        mem[946] = 32'b00111111111111110011111111111111;
        mem[947] = 32'b00111111111111110011111111111111;
        mem[948] = 32'b00111111111111110011111111111111;
        mem[949] = 32'b00111111111111110011111111111111;
        mem[950] = 32'b00111111111111110011111111111111;
        mem[951] = 32'b00111111111111110011111111111111;
        mem[952] = 32'b00111111111111110011111111111111;
        mem[953] = 32'b00111111111111110011111111111111;
        mem[954] = 32'b00111111111111110011111111111111;
        mem[955] = 32'b00111111111111110011111111111111;
        mem[956] = 32'b00111111111111110011111111111111;
        mem[957] = 32'b00111111111111110011111111111111;
        mem[958] = 32'b00111111111111110011111111111111;
        mem[959] = 32'b00111111111111110011111111111111;
        mem[960] = 32'b00111111111111110011111111111111;
        mem[961] = 32'b00111111111111110011111111111111;
        mem[962] = 32'b00111111111111110011111111111111;
        mem[963] = 32'b00111111111111110011111111111111;
        mem[964] = 32'b00111111111111110011111111111111;
        mem[965] = 32'b00111111111111110011111111111111;
        mem[966] = 32'b00111111111111110011111111111111;
        mem[967] = 32'b00111111111111110011111111111111;
        mem[968] = 32'b00111111111111110011111111111111;
        mem[969] = 32'b00111111111111110011111111111111;
        mem[970] = 32'b00111111111111110011111111111111;
        mem[971] = 32'b00111111111111110011111111111111;
        mem[972] = 32'b00111111111111110011111111111111;
        mem[973] = 32'b00111111111111110011111111111111;
        mem[974] = 32'b00111111111111110011111111111111;
        mem[975] = 32'b00111111111111110011111111111111;
        mem[976] = 32'b00111111111111110011111111111111;
        mem[977] = 32'b00111111111111110011111111111111;
        mem[978] = 32'b00111111111111110011111111111111;
        mem[979] = 32'b00111111111111110011111111111111;
        mem[980] = 32'b00111111111111110011111111111111;
        mem[981] = 32'b00111111111111110011111111111111;
        mem[982] = 32'b00111111111111110011111111111111;
        mem[983] = 32'b00111111111111110011111111111111;
        mem[984] = 32'b00111111111111110011111111111111;
        mem[985] = 32'b00111111111111110011111111111111;
        mem[986] = 32'b00111111111111110011111111111111;
        mem[987] = 32'b00111111111111110011111111111111;
        mem[988] = 32'b00111111111111110011111111111111;
        mem[989] = 32'b00111111111111110011111111111111;
        mem[990] = 32'b00111111111111110011111111111111;
        mem[991] = 32'b00111111111111110011111111111111;
        mem[992] = 32'b00111111111111110011111111111111;
        mem[993] = 32'b00111111111111110011111111111111;
        mem[994] = 32'b00111111111111110011111111111111;
        mem[995] = 32'b00111111111111110011111111111111;
        mem[996] = 32'b00111111111111110011111111111111;
        mem[997] = 32'b00111111111111110011111111111111;
        mem[998] = 32'b00111111111111110011111111111111;
        mem[999] = 32'b00111111111111110011111111111111;
        mem[1000] = 32'b00111111111111110011111111111111;
        mem[1001] = 32'b00111111111111110011111111111111;
        mem[1002] = 32'b00111111111111110011111111111111;
        mem[1003] = 32'b00111111111111110011111111111111;
        mem[1004] = 32'b00111111111111110011111111111111;
        mem[1005] = 32'b00111111111111110011111111111111;
        mem[1006] = 32'b00111111111111110011111111111111;
        mem[1007] = 32'b00111111111111110011111111111111;
        mem[1008] = 32'b00111111111111110011111111111111;
        mem[1009] = 32'b00111111111111110011111111111111;
        mem[1010] = 32'b00111111111111110011111111111111;
        mem[1011] = 32'b00111111111111110011111111111111;
        mem[1012] = 32'b00111111111111110011111111111111;
        mem[1013] = 32'b00111111111111110011111111111111;
        mem[1014] = 32'b00111111111111110011111111111111;
        mem[1015] = 32'b00111111111111110011111111111111;
        mem[1016] = 32'b00111111111111110011111111111111;
        mem[1017] = 32'b00111111111111110011111111111111;
        mem[1018] = 32'b00111111111111110011111111111111;
        mem[1019] = 32'b00111111111111110011111111111111;
        mem[1020] = 32'b00111111111111110011111111111111;
        mem[1021] = 32'b00111111111111110011111111111111;
        mem[1022] = 32'b00111111111111110011111111111111;
    end
endmodule