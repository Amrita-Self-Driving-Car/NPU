//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.08.2021 22:17:08
// Design Name: 
// Module Name: X_Rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module X_Rom(
  input load_mem
);
    reg [15:0] mem [1023:0];
    always @(posedge load_mem)
    begin
        mem[0] = 16'b1000000001000000;
        mem[1] = 16'b1000000010000000;
        mem[2] = 16'b1000000011000000;
        mem[3] = 16'b1000000100000000;
        mem[4] = 16'b1000000101000000;
        mem[5] = 16'b1000000110000000;
        mem[6] = 16'b1000000111000000;
        mem[7] = 16'b1000001000000000;
        mem[8] = 16'b1000001001000000;
        mem[9] = 16'b1000001010000000;
        mem[10] = 16'b1000001011000000;
        mem[11] = 16'b1000001100000000;
        mem[12] = 16'b1000001101000000;
        mem[13] = 16'b1000001110000000;
        mem[14] = 16'b1000001111000000;
        mem[15] = 16'b1000010000000000;
        mem[16] = 16'b1000010001000000;
        mem[17] = 16'b1000010010000000;
        mem[18] = 16'b1000010011000000;
        mem[19] = 16'b1000010100000000;
        mem[20] = 16'b1000010101000000;
        mem[21] = 16'b1000010110000000;
        mem[22] = 16'b1000010111000000;
        mem[23] = 16'b1000011000000000;
        mem[24] = 16'b1000011001000000;
        mem[25] = 16'b1000011010000000;
        mem[26] = 16'b1000011011000000;
        mem[27] = 16'b1000011100000000;
        mem[28] = 16'b1000011101000000;
        mem[29] = 16'b1000011110000000;
        mem[30] = 16'b1000011111000000;
        mem[31] = 16'b1000100000000000;
        mem[32] = 16'b1000100001000000;
        mem[33] = 16'b1000100010000000;
        mem[34] = 16'b1000100011000000;
        mem[35] = 16'b1000100100000000;
        mem[36] = 16'b1000100101000000;
        mem[37] = 16'b1000100110000000;
        mem[38] = 16'b1000100111000000;
        mem[39] = 16'b1000101000000000;
        mem[40] = 16'b1000101001000000;
        mem[41] = 16'b1000101010000000;
        mem[42] = 16'b1000101011000000;
        mem[43] = 16'b1000101100000000;
        mem[44] = 16'b1000101101000000;
        mem[45] = 16'b1000101110000000;
        mem[46] = 16'b1000101111000000;
        mem[47] = 16'b1000110000000000;
        mem[48] = 16'b1000110001000000;
        mem[49] = 16'b1000110010000000;
        mem[50] = 16'b1000110011000000;
        mem[51] = 16'b1000110100000000;
        mem[52] = 16'b1000110101000000;
        mem[53] = 16'b1000110110000000;
        mem[54] = 16'b1000110111000000;
        mem[55] = 16'b1000111000000000;
        mem[56] = 16'b1000111001000000;
        mem[57] = 16'b1000111010000000;
        mem[58] = 16'b1000111011000000;
        mem[59] = 16'b1000111100000000;
        mem[60] = 16'b1000111101000000;
        mem[61] = 16'b1000111110000000;
        mem[62] = 16'b1000111111000000;
        mem[63] = 16'b1001000000000000;
        mem[64] = 16'b1001000001000000;
        mem[65] = 16'b1001000010000000;
        mem[66] = 16'b1001000011000000;
        mem[67] = 16'b1001000100000000;
        mem[68] = 16'b1001000101000000;
        mem[69] = 16'b1001000110000000;
        mem[70] = 16'b1001000111000000;
        mem[71] = 16'b1001001000000000;
        mem[72] = 16'b1001001001000000;
        mem[73] = 16'b1001001010000000;
        mem[74] = 16'b1001001011000000;
        mem[75] = 16'b1001001100000000;
        mem[76] = 16'b1001001101000000;
        mem[77] = 16'b1001001110000000;
        mem[78] = 16'b1001001111000000;
        mem[79] = 16'b1001010000000000;
        mem[80] = 16'b1001010001000000;
        mem[81] = 16'b1001010010000000;
        mem[82] = 16'b1001010011000000;
        mem[83] = 16'b1001010100000000;
        mem[84] = 16'b1001010101000000;
        mem[85] = 16'b1001010110000000;
        mem[86] = 16'b1001010111000000;
        mem[87] = 16'b1001011000000000;
        mem[88] = 16'b1001011001000000;
        mem[89] = 16'b1001011010000000;
        mem[90] = 16'b1001011011000000;
        mem[91] = 16'b1001011100000000;
        mem[92] = 16'b1001011101000000;
        mem[93] = 16'b1001011110000000;
        mem[94] = 16'b1001011111000000;
        mem[95] = 16'b1001100000000000;
        mem[96] = 16'b1001100001000000;
        mem[97] = 16'b1001100010000000;
        mem[98] = 16'b1001100011000000;
        mem[99] = 16'b1001100100000000;
        mem[100] = 16'b1001100101000000;
        mem[101] = 16'b1001100110000000;
        mem[102] = 16'b1001100111000000;
        mem[103] = 16'b1001101000000000;
        mem[104] = 16'b1001101001000000;
        mem[105] = 16'b1001101010000000;
        mem[106] = 16'b1001101011000000;
        mem[107] = 16'b1001101100000000;
        mem[108] = 16'b1001101101000000;
        mem[109] = 16'b1001101110000000;
        mem[110] = 16'b1001101111000000;
        mem[111] = 16'b1001110000000000;
        mem[112] = 16'b1001110001000000;
        mem[113] = 16'b1001110010000000;
        mem[114] = 16'b1001110011000000;
        mem[115] = 16'b1001110100000000;
        mem[116] = 16'b1001110101000000;
        mem[117] = 16'b1001110110000000;
        mem[118] = 16'b1001110111000000;
        mem[119] = 16'b1001111000000000;
        mem[120] = 16'b1001111001000000;
        mem[121] = 16'b1001111010000000;
        mem[122] = 16'b1001111011000000;
        mem[123] = 16'b1001111100000000;
        mem[124] = 16'b1001111101000000;
        mem[125] = 16'b1001111110000000;
        mem[126] = 16'b1001111111000000;
        mem[127] = 16'b1010000000000000;
        mem[128] = 16'b1010000001000000;
        mem[129] = 16'b1010000010000000;
        mem[130] = 16'b1010000011000000;
        mem[131] = 16'b1010000100000000;
        mem[132] = 16'b1010000101000000;
        mem[133] = 16'b1010000110000000;
        mem[134] = 16'b1010000111000000;
        mem[135] = 16'b1010001000000000;
        mem[136] = 16'b1010001001000000;
        mem[137] = 16'b1010001010000000;
        mem[138] = 16'b1010001011000000;
        mem[139] = 16'b1010001100000000;
        mem[140] = 16'b1010001101000000;
        mem[141] = 16'b1010001110000000;
        mem[142] = 16'b1010001111000000;
        mem[143] = 16'b1010010000000000;
        mem[144] = 16'b1010010001000000;
        mem[145] = 16'b1010010010000000;
        mem[146] = 16'b1010010011000000;
        mem[147] = 16'b1010010100000000;
        mem[148] = 16'b1010010101000000;
        mem[149] = 16'b1010010110000000;
        mem[150] = 16'b1010010111000000;
        mem[151] = 16'b1010011000000000;
        mem[152] = 16'b1010011001000000;
        mem[153] = 16'b1010011010000000;
        mem[154] = 16'b1010011011000000;
        mem[155] = 16'b1010011100000000;
        mem[156] = 16'b1010011101000000;
        mem[157] = 16'b1010011110000000;
        mem[158] = 16'b1010011111000000;
        mem[159] = 16'b1010100000000000;
        mem[160] = 16'b1010100001000000;
        mem[161] = 16'b1010100010000000;
        mem[162] = 16'b1010100011000000;
        mem[163] = 16'b1010100100000000;
        mem[164] = 16'b1010100101000000;
        mem[165] = 16'b1010100110000000;
        mem[166] = 16'b1010100111000000;
        mem[167] = 16'b1010101000000000;
        mem[168] = 16'b1010101001000000;
        mem[169] = 16'b1010101010000000;
        mem[170] = 16'b1010101011000000;
        mem[171] = 16'b1010101100000000;
        mem[172] = 16'b1010101101000000;
        mem[173] = 16'b1010101110000000;
        mem[174] = 16'b1010101111000000;
        mem[175] = 16'b1010110000000000;
        mem[176] = 16'b1010110001000000;
        mem[177] = 16'b1010110010000000;
        mem[178] = 16'b1010110011000000;
        mem[179] = 16'b1010110100000000;
        mem[180] = 16'b1010110101000000;
        mem[181] = 16'b1010110110000000;
        mem[182] = 16'b1010110111000000;
        mem[183] = 16'b1010111000000000;
        mem[184] = 16'b1010111001000000;
        mem[185] = 16'b1010111010000000;
        mem[186] = 16'b1010111011000000;
        mem[187] = 16'b1010111100000000;
        mem[188] = 16'b1010111101000000;
        mem[189] = 16'b1010111110000000;
        mem[190] = 16'b1010111111000000;
        mem[191] = 16'b1011000000000000;
        mem[192] = 16'b1011000001000000;
        mem[193] = 16'b1011000010000000;
        mem[194] = 16'b1011000011000000;
        mem[195] = 16'b1011000100000000;
        mem[196] = 16'b1011000101000000;
        mem[197] = 16'b1011000110000000;
        mem[198] = 16'b1011000111000000;
        mem[199] = 16'b1011001000000000;
        mem[200] = 16'b1011001001000000;
        mem[201] = 16'b1011001010000000;
        mem[202] = 16'b1011001011000000;
        mem[203] = 16'b1011001100000000;
        mem[204] = 16'b1011001101000000;
        mem[205] = 16'b1011001110000000;
        mem[206] = 16'b1011001111000000;
        mem[207] = 16'b1011010000000000;
        mem[208] = 16'b1011010001000000;
        mem[209] = 16'b1011010010000000;
        mem[210] = 16'b1011010011000000;
        mem[211] = 16'b1011010100000000;
        mem[212] = 16'b1011010101000000;
        mem[213] = 16'b1011010110000000;
        mem[214] = 16'b1011010111000000;
        mem[215] = 16'b1011011000000000;
        mem[216] = 16'b1011011001000000;
        mem[217] = 16'b1011011010000000;
        mem[218] = 16'b1011011011000000;
        mem[219] = 16'b1011011100000000;
        mem[220] = 16'b1011011101000000;
        mem[221] = 16'b1011011110000000;
        mem[222] = 16'b1011011111000000;
        mem[223] = 16'b1011100000000000;
        mem[224] = 16'b1011100001000000;
        mem[225] = 16'b1011100010000000;
        mem[226] = 16'b1011100011000000;
        mem[227] = 16'b1011100100000000;
        mem[228] = 16'b1011100101000000;
        mem[229] = 16'b1011100110000000;
        mem[230] = 16'b1011100111000000;
        mem[231] = 16'b1011101000000000;
        mem[232] = 16'b1011101001000000;
        mem[233] = 16'b1011101010000000;
        mem[234] = 16'b1011101011000000;
        mem[235] = 16'b1011101100000000;
        mem[236] = 16'b1011101101000000;
        mem[237] = 16'b1011101110000000;
        mem[238] = 16'b1011101111000000;
        mem[239] = 16'b1011110000000000;
        mem[240] = 16'b1011110001000000;
        mem[241] = 16'b1011110010000000;
        mem[242] = 16'b1011110011000000;
        mem[243] = 16'b1011110100000000;
        mem[244] = 16'b1011110101000000;
        mem[245] = 16'b1011110110000000;
        mem[246] = 16'b1011110111000000;
        mem[247] = 16'b1011111000000000;
        mem[248] = 16'b1011111001000000;
        mem[249] = 16'b1011111010000000;
        mem[250] = 16'b1011111011000000;
        mem[251] = 16'b1011111100000000;
        mem[252] = 16'b1011111101000000;
        mem[253] = 16'b1011111110000000;
        mem[254] = 16'b1011111111000000;
        mem[255] = 16'b1100000000000000;
        mem[256] = 16'b1100000001000000;
        mem[257] = 16'b1100000010000000;
        mem[258] = 16'b1100000011000000;
        mem[259] = 16'b1100000100000000;
        mem[260] = 16'b1100000101000000;
        mem[261] = 16'b1100000110000000;
        mem[262] = 16'b1100000111000000;
        mem[263] = 16'b1100001000000000;
        mem[264] = 16'b1100001001000000;
        mem[265] = 16'b1100001010000000;
        mem[266] = 16'b1100001011000000;
        mem[267] = 16'b1100001100000000;
        mem[268] = 16'b1100001101000000;
        mem[269] = 16'b1100001110000000;
        mem[270] = 16'b1100001111000000;
        mem[271] = 16'b1100010000000000;
        mem[272] = 16'b1100010001000000;
        mem[273] = 16'b1100010010000000;
        mem[274] = 16'b1100010011000000;
        mem[275] = 16'b1100010100000000;
        mem[276] = 16'b1100010101000000;
        mem[277] = 16'b1100010110000000;
        mem[278] = 16'b1100010111000000;
        mem[279] = 16'b1100011000000000;
        mem[280] = 16'b1100011001000000;
        mem[281] = 16'b1100011010000000;
        mem[282] = 16'b1100011011000000;
        mem[283] = 16'b1100011100000000;
        mem[284] = 16'b1100011101000000;
        mem[285] = 16'b1100011110000000;
        mem[286] = 16'b1100011111000000;
        mem[287] = 16'b1100100000000000;
        mem[288] = 16'b1100100001000000;
        mem[289] = 16'b1100100010000000;
        mem[290] = 16'b1100100011000000;
        mem[291] = 16'b1100100100000000;
        mem[292] = 16'b1100100101000000;
        mem[293] = 16'b1100100110000000;
        mem[294] = 16'b1100100111000000;
        mem[295] = 16'b1100101000000000;
        mem[296] = 16'b1100101001000000;
        mem[297] = 16'b1100101010000000;
        mem[298] = 16'b1100101011000000;
        mem[299] = 16'b1100101100000000;
        mem[300] = 16'b1100101101000000;
        mem[301] = 16'b1100101110000000;
        mem[302] = 16'b1100101111000000;
        mem[303] = 16'b1100110000000000;
        mem[304] = 16'b1100110001000000;
        mem[305] = 16'b1100110010000000;
        mem[306] = 16'b1100110011000000;
        mem[307] = 16'b1100110100000000;
        mem[308] = 16'b1100110101000000;
        mem[309] = 16'b1100110110000000;
        mem[310] = 16'b1100110111000000;
        mem[311] = 16'b1100111000000000;
        mem[312] = 16'b1100111001000000;
        mem[313] = 16'b1100111010000000;
        mem[314] = 16'b1100111011000000;
        mem[315] = 16'b1100111100000000;
        mem[316] = 16'b1100111101000000;
        mem[317] = 16'b1100111110000000;
        mem[318] = 16'b1100111111000000;
        mem[319] = 16'b1101000000000000;
        mem[320] = 16'b1101000001000000;
        mem[321] = 16'b1101000010000000;
        mem[322] = 16'b1101000011000000;
        mem[323] = 16'b1101000100000000;
        mem[324] = 16'b1101000101000000;
        mem[325] = 16'b1101000110000000;
        mem[326] = 16'b1101000111000000;
        mem[327] = 16'b1101001000000000;
        mem[328] = 16'b1101001001000000;
        mem[329] = 16'b1101001010000000;
        mem[330] = 16'b1101001011000000;
        mem[331] = 16'b1101001100000000;
        mem[332] = 16'b1101001101000000;
        mem[333] = 16'b1101001110000000;
        mem[334] = 16'b1101001111000000;
        mem[335] = 16'b1101010000000000;
        mem[336] = 16'b1101010001000000;
        mem[337] = 16'b1101010010000000;
        mem[338] = 16'b1101010011000000;
        mem[339] = 16'b1101010100000000;
        mem[340] = 16'b1101010101000000;
        mem[341] = 16'b1101010110000000;
        mem[342] = 16'b1101010111000000;
        mem[343] = 16'b1101011000000000;
        mem[344] = 16'b1101011001000000;
        mem[345] = 16'b1101011010000000;
        mem[346] = 16'b1101011011000000;
        mem[347] = 16'b1101011100000000;
        mem[348] = 16'b1101011101000000;
        mem[349] = 16'b1101011110000000;
        mem[350] = 16'b1101011111000000;
        mem[351] = 16'b1101100000000000;
        mem[352] = 16'b1101100001000000;
        mem[353] = 16'b1101100010000000;
        mem[354] = 16'b1101100011000000;
        mem[355] = 16'b1101100100000000;
        mem[356] = 16'b1101100101000000;
        mem[357] = 16'b1101100110000000;
        mem[358] = 16'b1101100111000000;
        mem[359] = 16'b1101101000000000;
        mem[360] = 16'b1101101001000000;
        mem[361] = 16'b1101101010000000;
        mem[362] = 16'b1101101011000000;
        mem[363] = 16'b1101101100000000;
        mem[364] = 16'b1101101101000000;
        mem[365] = 16'b1101101110000000;
        mem[366] = 16'b1101101111000000;
        mem[367] = 16'b1101110000000000;
        mem[368] = 16'b1101110001000000;
        mem[369] = 16'b1101110010000000;
        mem[370] = 16'b1101110011000000;
        mem[371] = 16'b1101110100000000;
        mem[372] = 16'b1101110101000000;
        mem[373] = 16'b1101110110000000;
        mem[374] = 16'b1101110111000000;
        mem[375] = 16'b1101111000000000;
        mem[376] = 16'b1101111001000000;
        mem[377] = 16'b1101111010000000;
        mem[378] = 16'b1101111011000000;
        mem[379] = 16'b1101111100000000;
        mem[380] = 16'b1101111101000000;
        mem[381] = 16'b1101111110000000;
        mem[382] = 16'b1101111111000000;
        mem[383] = 16'b1110000000000000;
        mem[384] = 16'b1110000001000000;
        mem[385] = 16'b1110000010000000;
        mem[386] = 16'b1110000011000000;
        mem[387] = 16'b1110000100000000;
        mem[388] = 16'b1110000101000000;
        mem[389] = 16'b1110000110000000;
        mem[390] = 16'b1110000111000000;
        mem[391] = 16'b1110001000000000;
        mem[392] = 16'b1110001001000000;
        mem[393] = 16'b1110001010000000;
        mem[394] = 16'b1110001011000000;
        mem[395] = 16'b1110001100000000;
        mem[396] = 16'b1110001101000000;
        mem[397] = 16'b1110001110000000;
        mem[398] = 16'b1110001111000000;
        mem[399] = 16'b1110010000000000;
        mem[400] = 16'b1110010001000000;
        mem[401] = 16'b1110010010000000;
        mem[402] = 16'b1110010011000000;
        mem[403] = 16'b1110010100000000;
        mem[404] = 16'b1110010101000000;
        mem[405] = 16'b1110010110000000;
        mem[406] = 16'b1110010111000000;
        mem[407] = 16'b1110011000000000;
        mem[408] = 16'b1110011001000000;
        mem[409] = 16'b1110011010000000;
        mem[410] = 16'b1110011011000000;
        mem[411] = 16'b1110011100000000;
        mem[412] = 16'b1110011101000000;
        mem[413] = 16'b1110011110000000;
        mem[414] = 16'b1110011111000000;
        mem[415] = 16'b1110100000000000;
        mem[416] = 16'b1110100001000000;
        mem[417] = 16'b1110100010000000;
        mem[418] = 16'b1110100011000000;
        mem[419] = 16'b1110100100000000;
        mem[420] = 16'b1110100101000000;
        mem[421] = 16'b1110100110000000;
        mem[422] = 16'b1110100111000000;
        mem[423] = 16'b1110101000000000;
        mem[424] = 16'b1110101001000000;
        mem[425] = 16'b1110101010000000;
        mem[426] = 16'b1110101011000000;
        mem[427] = 16'b1110101100000000;
        mem[428] = 16'b1110101101000000;
        mem[429] = 16'b1110101110000000;
        mem[430] = 16'b1110101111000000;
        mem[431] = 16'b1110110000000000;
        mem[432] = 16'b1110110001000000;
        mem[433] = 16'b1110110010000000;
        mem[434] = 16'b1110110011000000;
        mem[435] = 16'b1110110100000000;
        mem[436] = 16'b1110110101000000;
        mem[437] = 16'b1110110110000000;
        mem[438] = 16'b1110110111000000;
        mem[439] = 16'b1110111000000000;
        mem[440] = 16'b1110111001000000;
        mem[441] = 16'b1110111010000000;
        mem[442] = 16'b1110111011000000;
        mem[443] = 16'b1110111100000000;
        mem[444] = 16'b1110111101000000;
        mem[445] = 16'b1110111110000000;
        mem[446] = 16'b1110111111000000;
        mem[447] = 16'b1111000000000000;
        mem[448] = 16'b1111000001000000;
        mem[449] = 16'b1111000010000000;
        mem[450] = 16'b1111000011000000;
        mem[451] = 16'b1111000100000000;
        mem[452] = 16'b1111000101000000;
        mem[453] = 16'b1111000110000000;
        mem[454] = 16'b1111000111000000;
        mem[455] = 16'b1111001000000000;
        mem[456] = 16'b1111001001000000;
        mem[457] = 16'b1111001010000000;
        mem[458] = 16'b1111001011000000;
        mem[459] = 16'b1111001100000000;
        mem[460] = 16'b1111001101000000;
        mem[461] = 16'b1111001110000000;
        mem[462] = 16'b1111001111000000;
        mem[463] = 16'b1111010000000000;
        mem[464] = 16'b1111010001000000;
        mem[465] = 16'b1111010010000000;
        mem[466] = 16'b1111010011000000;
        mem[467] = 16'b1111010100000000;
        mem[468] = 16'b1111010101000000;
        mem[469] = 16'b1111010110000000;
        mem[470] = 16'b1111010111000000;
        mem[471] = 16'b1111011000000000;
        mem[472] = 16'b1111011001000000;
        mem[473] = 16'b1111011010000000;
        mem[474] = 16'b1111011011000000;
        mem[475] = 16'b1111011100000000;
        mem[476] = 16'b1111011101000000;
        mem[477] = 16'b1111011110000000;
        mem[478] = 16'b1111011111000000;
        mem[479] = 16'b1111100000000000;
        mem[480] = 16'b1111100001000000;
        mem[481] = 16'b1111100010000000;
        mem[482] = 16'b1111100011000000;
        mem[483] = 16'b1111100100000000;
        mem[484] = 16'b1111100101000000;
        mem[485] = 16'b1111100110000000;
        mem[486] = 16'b1111100111000000;
        mem[487] = 16'b1111101000000000;
        mem[488] = 16'b1111101001000000;
        mem[489] = 16'b1111101010000000;
        mem[490] = 16'b1111101011000000;
        mem[491] = 16'b1111101100000000;
        mem[492] = 16'b1111101101000000;
        mem[493] = 16'b1111101110000000;
        mem[494] = 16'b1111101111000000;
        mem[495] = 16'b1111110000000000;
        mem[496] = 16'b1111110001000000;
        mem[497] = 16'b1111110010000000;
        mem[498] = 16'b1111110011000000;
        mem[499] = 16'b1111110100000000;
        mem[500] = 16'b1111110101000000;
        mem[501] = 16'b1111110110000000;
        mem[502] = 16'b1111110111000000;
        mem[503] = 16'b1111111000000000;
        mem[504] = 16'b1111111001000000;
        mem[505] = 16'b1111111010000000;
        mem[506] = 16'b1111111011000000;
        mem[507] = 16'b1111111100000000;
        mem[508] = 16'b1111111101000000;
        mem[509] = 16'b1111111110000000;
        mem[510] = 16'b1111111111000000;
        mem[511] = 16'b0000000000000000;
        mem[512] = 16'b0000000001000000;
        mem[513] = 16'b0000000010000000;
        mem[514] = 16'b0000000011000000;
        mem[515] = 16'b0000000100000000;
        mem[516] = 16'b0000000101000000;
        mem[517] = 16'b0000000110000000;
        mem[518] = 16'b0000000111000000;
        mem[519] = 16'b0000001000000000;
        mem[520] = 16'b0000001001000000;
        mem[521] = 16'b0000001010000000;
        mem[522] = 16'b0000001011000000;
        mem[523] = 16'b0000001100000000;
        mem[524] = 16'b0000001101000000;
        mem[525] = 16'b0000001110000000;
        mem[526] = 16'b0000001111000000;
        mem[527] = 16'b0000010000000000;
        mem[528] = 16'b0000010001000000;
        mem[529] = 16'b0000010010000000;
        mem[530] = 16'b0000010011000000;
        mem[531] = 16'b0000010100000000;
        mem[532] = 16'b0000010101000000;
        mem[533] = 16'b0000010110000000;
        mem[534] = 16'b0000010111000000;
        mem[535] = 16'b0000011000000000;
        mem[536] = 16'b0000011001000000;
        mem[537] = 16'b0000011010000000;
        mem[538] = 16'b0000011011000000;
        mem[539] = 16'b0000011100000000;
        mem[540] = 16'b0000011101000000;
        mem[541] = 16'b0000011110000000;
        mem[542] = 16'b0000011111000000;
        mem[543] = 16'b0000100000000000;
        mem[544] = 16'b0000100001000000;
        mem[545] = 16'b0000100010000000;
        mem[546] = 16'b0000100011000000;
        mem[547] = 16'b0000100100000000;
        mem[548] = 16'b0000100101000000;
        mem[549] = 16'b0000100110000000;
        mem[550] = 16'b0000100111000000;
        mem[551] = 16'b0000101000000000;
        mem[552] = 16'b0000101001000000;
        mem[553] = 16'b0000101010000000;
        mem[554] = 16'b0000101011000000;
        mem[555] = 16'b0000101100000000;
        mem[556] = 16'b0000101101000000;
        mem[557] = 16'b0000101110000000;
        mem[558] = 16'b0000101111000000;
        mem[559] = 16'b0000110000000000;
        mem[560] = 16'b0000110001000000;
        mem[561] = 16'b0000110010000000;
        mem[562] = 16'b0000110011000000;
        mem[563] = 16'b0000110100000000;
        mem[564] = 16'b0000110101000000;
        mem[565] = 16'b0000110110000000;
        mem[566] = 16'b0000110111000000;
        mem[567] = 16'b0000111000000000;
        mem[568] = 16'b0000111001000000;
        mem[569] = 16'b0000111010000000;
        mem[570] = 16'b0000111011000000;
        mem[571] = 16'b0000111100000000;
        mem[572] = 16'b0000111101000000;
        mem[573] = 16'b0000111110000000;
        mem[574] = 16'b0000111111000000;
        mem[575] = 16'b0001000000000000;
        mem[576] = 16'b0001000001000000;
        mem[577] = 16'b0001000010000000;
        mem[578] = 16'b0001000011000000;
        mem[579] = 16'b0001000100000000;
        mem[580] = 16'b0001000101000000;
        mem[581] = 16'b0001000110000000;
        mem[582] = 16'b0001000111000000;
        mem[583] = 16'b0001001000000000;
        mem[584] = 16'b0001001001000000;
        mem[585] = 16'b0001001010000000;
        mem[586] = 16'b0001001011000000;
        mem[587] = 16'b0001001100000000;
        mem[588] = 16'b0001001101000000;
        mem[589] = 16'b0001001110000000;
        mem[590] = 16'b0001001111000000;
        mem[591] = 16'b0001010000000000;
        mem[592] = 16'b0001010001000000;
        mem[593] = 16'b0001010010000000;
        mem[594] = 16'b0001010011000000;
        mem[595] = 16'b0001010100000000;
        mem[596] = 16'b0001010101000000;
        mem[597] = 16'b0001010110000000;
        mem[598] = 16'b0001010111000000;
        mem[599] = 16'b0001011000000000;
        mem[600] = 16'b0001011001000000;
        mem[601] = 16'b0001011010000000;
        mem[602] = 16'b0001011011000000;
        mem[603] = 16'b0001011100000000;
        mem[604] = 16'b0001011101000000;
        mem[605] = 16'b0001011110000000;
        mem[606] = 16'b0001011111000000;
        mem[607] = 16'b0001100000000000;
        mem[608] = 16'b0001100001000000;
        mem[609] = 16'b0001100010000000;
        mem[610] = 16'b0001100011000000;
        mem[611] = 16'b0001100100000000;
        mem[612] = 16'b0001100101000000;
        mem[613] = 16'b0001100110000000;
        mem[614] = 16'b0001100111000000;
        mem[615] = 16'b0001101000000000;
        mem[616] = 16'b0001101001000000;
        mem[617] = 16'b0001101010000000;
        mem[618] = 16'b0001101011000000;
        mem[619] = 16'b0001101100000000;
        mem[620] = 16'b0001101101000000;
        mem[621] = 16'b0001101110000000;
        mem[622] = 16'b0001101111000000;
        mem[623] = 16'b0001110000000000;
        mem[624] = 16'b0001110001000000;
        mem[625] = 16'b0001110010000000;
        mem[626] = 16'b0001110011000000;
        mem[627] = 16'b0001110100000000;
        mem[628] = 16'b0001110101000000;
        mem[629] = 16'b0001110110000000;
        mem[630] = 16'b0001110111000000;
        mem[631] = 16'b0001111000000000;
        mem[632] = 16'b0001111001000000;
        mem[633] = 16'b0001111010000000;
        mem[634] = 16'b0001111011000000;
        mem[635] = 16'b0001111100000000;
        mem[636] = 16'b0001111101000000;
        mem[637] = 16'b0001111110000000;
        mem[638] = 16'b0001111111000000;
        mem[639] = 16'b0010000000000000;
        mem[640] = 16'b0010000001000000;
        mem[641] = 16'b0010000010000000;
        mem[642] = 16'b0010000011000000;
        mem[643] = 16'b0010000100000000;
        mem[644] = 16'b0010000101000000;
        mem[645] = 16'b0010000110000000;
        mem[646] = 16'b0010000111000000;
        mem[647] = 16'b0010001000000000;
        mem[648] = 16'b0010001001000000;
        mem[649] = 16'b0010001010000000;
        mem[650] = 16'b0010001011000000;
        mem[651] = 16'b0010001100000000;
        mem[652] = 16'b0010001101000000;
        mem[653] = 16'b0010001110000000;
        mem[654] = 16'b0010001111000000;
        mem[655] = 16'b0010010000000000;
        mem[656] = 16'b0010010001000000;
        mem[657] = 16'b0010010010000000;
        mem[658] = 16'b0010010011000000;
        mem[659] = 16'b0010010100000000;
        mem[660] = 16'b0010010101000000;
        mem[661] = 16'b0010010110000000;
        mem[662] = 16'b0010010111000000;
        mem[663] = 16'b0010011000000000;
        mem[664] = 16'b0010011001000000;
        mem[665] = 16'b0010011010000000;
        mem[666] = 16'b0010011011000000;
        mem[667] = 16'b0010011100000000;
        mem[668] = 16'b0010011101000000;
        mem[669] = 16'b0010011110000000;
        mem[670] = 16'b0010011111000000;
        mem[671] = 16'b0010100000000000;
        mem[672] = 16'b0010100001000000;
        mem[673] = 16'b0010100010000000;
        mem[674] = 16'b0010100011000000;
        mem[675] = 16'b0010100100000000;
        mem[676] = 16'b0010100101000000;
        mem[677] = 16'b0010100110000000;
        mem[678] = 16'b0010100111000000;
        mem[679] = 16'b0010101000000000;
        mem[680] = 16'b0010101001000000;
        mem[681] = 16'b0010101010000000;
        mem[682] = 16'b0010101011000000;
        mem[683] = 16'b0010101100000000;
        mem[684] = 16'b0010101101000000;
        mem[685] = 16'b0010101110000000;
        mem[686] = 16'b0010101111000000;
        mem[687] = 16'b0010110000000000;
        mem[688] = 16'b0010110001000000;
        mem[689] = 16'b0010110010000000;
        mem[690] = 16'b0010110011000000;
        mem[691] = 16'b0010110100000000;
        mem[692] = 16'b0010110101000000;
        mem[693] = 16'b0010110110000000;
        mem[694] = 16'b0010110111000000;
        mem[695] = 16'b0010111000000000;
        mem[696] = 16'b0010111001000000;
        mem[697] = 16'b0010111010000000;
        mem[698] = 16'b0010111011000000;
        mem[699] = 16'b0010111100000000;
        mem[700] = 16'b0010111101000000;
        mem[701] = 16'b0010111110000000;
        mem[702] = 16'b0010111111000000;
        mem[703] = 16'b0011000000000000;
        mem[704] = 16'b0011000001000000;
        mem[705] = 16'b0011000010000000;
        mem[706] = 16'b0011000011000000;
        mem[707] = 16'b0011000100000000;
        mem[708] = 16'b0011000101000000;
        mem[709] = 16'b0011000110000000;
        mem[710] = 16'b0011000111000000;
        mem[711] = 16'b0011001000000000;
        mem[712] = 16'b0011001001000000;
        mem[713] = 16'b0011001010000000;
        mem[714] = 16'b0011001011000000;
        mem[715] = 16'b0011001100000000;
        mem[716] = 16'b0011001101000000;
        mem[717] = 16'b0011001110000000;
        mem[718] = 16'b0011001111000000;
        mem[719] = 16'b0011010000000000;
        mem[720] = 16'b0011010001000000;
        mem[721] = 16'b0011010010000000;
        mem[722] = 16'b0011010011000000;
        mem[723] = 16'b0011010100000000;
        mem[724] = 16'b0011010101000000;
        mem[725] = 16'b0011010110000000;
        mem[726] = 16'b0011010111000000;
        mem[727] = 16'b0011011000000000;
        mem[728] = 16'b0011011001000000;
        mem[729] = 16'b0011011010000000;
        mem[730] = 16'b0011011011000000;
        mem[731] = 16'b0011011100000000;
        mem[732] = 16'b0011011101000000;
        mem[733] = 16'b0011011110000000;
        mem[734] = 16'b0011011111000000;
        mem[735] = 16'b0011100000000000;
        mem[736] = 16'b0011100001000000;
        mem[737] = 16'b0011100010000000;
        mem[738] = 16'b0011100011000000;
        mem[739] = 16'b0011100100000000;
        mem[740] = 16'b0011100101000000;
        mem[741] = 16'b0011100110000000;
        mem[742] = 16'b0011100111000000;
        mem[743] = 16'b0011101000000000;
        mem[744] = 16'b0011101001000000;
        mem[745] = 16'b0011101010000000;
        mem[746] = 16'b0011101011000000;
        mem[747] = 16'b0011101100000000;
        mem[748] = 16'b0011101101000000;
        mem[749] = 16'b0011101110000000;
        mem[750] = 16'b0011101111000000;
        mem[751] = 16'b0011110000000000;
        mem[752] = 16'b0011110001000000;
        mem[753] = 16'b0011110010000000;
        mem[754] = 16'b0011110011000000;
        mem[755] = 16'b0011110100000000;
        mem[756] = 16'b0011110101000000;
        mem[757] = 16'b0011110110000000;
        mem[758] = 16'b0011110111000000;
        mem[759] = 16'b0011111000000000;
        mem[760] = 16'b0011111001000000;
        mem[761] = 16'b0011111010000000;
        mem[762] = 16'b0011111011000000;
        mem[763] = 16'b0011111100000000;
        mem[764] = 16'b0011111101000000;
        mem[765] = 16'b0011111110000000;
        mem[766] = 16'b0011111111000000;
        mem[767] = 16'b0100000000000000;
        mem[768] = 16'b0100000001000000;
        mem[769] = 16'b0100000010000000;
        mem[770] = 16'b0100000011000000;
        mem[771] = 16'b0100000100000000;
        mem[772] = 16'b0100000101000000;
        mem[773] = 16'b0100000110000000;
        mem[774] = 16'b0100000111000000;
        mem[775] = 16'b0100001000000000;
        mem[776] = 16'b0100001001000000;
        mem[777] = 16'b0100001010000000;
        mem[778] = 16'b0100001011000000;
        mem[779] = 16'b0100001100000000;
        mem[780] = 16'b0100001101000000;
        mem[781] = 16'b0100001110000000;
        mem[782] = 16'b0100001111000000;
        mem[783] = 16'b0100010000000000;
        mem[784] = 16'b0100010001000000;
        mem[785] = 16'b0100010010000000;
        mem[786] = 16'b0100010011000000;
        mem[787] = 16'b0100010100000000;
        mem[788] = 16'b0100010101000000;
        mem[789] = 16'b0100010110000000;
        mem[790] = 16'b0100010111000000;
        mem[791] = 16'b0100011000000000;
        mem[792] = 16'b0100011001000000;
        mem[793] = 16'b0100011010000000;
        mem[794] = 16'b0100011011000000;
        mem[795] = 16'b0100011100000000;
        mem[796] = 16'b0100011101000000;
        mem[797] = 16'b0100011110000000;
        mem[798] = 16'b0100011111000000;
        mem[799] = 16'b0100100000000000;
        mem[800] = 16'b0100100001000000;
        mem[801] = 16'b0100100010000000;
        mem[802] = 16'b0100100011000000;
        mem[803] = 16'b0100100100000000;
        mem[804] = 16'b0100100101000000;
        mem[805] = 16'b0100100110000000;
        mem[806] = 16'b0100100111000000;
        mem[807] = 16'b0100101000000000;
        mem[808] = 16'b0100101001000000;
        mem[809] = 16'b0100101010000000;
        mem[810] = 16'b0100101011000000;
        mem[811] = 16'b0100101100000000;
        mem[812] = 16'b0100101101000000;
        mem[813] = 16'b0100101110000000;
        mem[814] = 16'b0100101111000000;
        mem[815] = 16'b0100110000000000;
        mem[816] = 16'b0100110001000000;
        mem[817] = 16'b0100110010000000;
        mem[818] = 16'b0100110011000000;
        mem[819] = 16'b0100110100000000;
        mem[820] = 16'b0100110101000000;
        mem[821] = 16'b0100110110000000;
        mem[822] = 16'b0100110111000000;
        mem[823] = 16'b0100111000000000;
        mem[824] = 16'b0100111001000000;
        mem[825] = 16'b0100111010000000;
        mem[826] = 16'b0100111011000000;
        mem[827] = 16'b0100111100000000;
        mem[828] = 16'b0100111101000000;
        mem[829] = 16'b0100111110000000;
        mem[830] = 16'b0100111111000000;
        mem[831] = 16'b0101000000000000;
        mem[832] = 16'b0101000001000000;
        mem[833] = 16'b0101000010000000;
        mem[834] = 16'b0101000011000000;
        mem[835] = 16'b0101000100000000;
        mem[836] = 16'b0101000101000000;
        mem[837] = 16'b0101000110000000;
        mem[838] = 16'b0101000111000000;
        mem[839] = 16'b0101001000000000;
        mem[840] = 16'b0101001001000000;
        mem[841] = 16'b0101001010000000;
        mem[842] = 16'b0101001011000000;
        mem[843] = 16'b0101001100000000;
        mem[844] = 16'b0101001101000000;
        mem[845] = 16'b0101001110000000;
        mem[846] = 16'b0101001111000000;
        mem[847] = 16'b0101010000000000;
        mem[848] = 16'b0101010001000000;
        mem[849] = 16'b0101010010000000;
        mem[850] = 16'b0101010011000000;
        mem[851] = 16'b0101010100000000;
        mem[852] = 16'b0101010101000000;
        mem[853] = 16'b0101010110000000;
        mem[854] = 16'b0101010111000000;
        mem[855] = 16'b0101011000000000;
        mem[856] = 16'b0101011001000000;
        mem[857] = 16'b0101011010000000;
        mem[858] = 16'b0101011011000000;
        mem[859] = 16'b0101011100000000;
        mem[860] = 16'b0101011101000000;
        mem[861] = 16'b0101011110000000;
        mem[862] = 16'b0101011111000000;
        mem[863] = 16'b0101100000000000;
        mem[864] = 16'b0101100001000000;
        mem[865] = 16'b0101100010000000;
        mem[866] = 16'b0101100011000000;
        mem[867] = 16'b0101100100000000;
        mem[868] = 16'b0101100101000000;
        mem[869] = 16'b0101100110000000;
        mem[870] = 16'b0101100111000000;
        mem[871] = 16'b0101101000000000;
        mem[872] = 16'b0101101001000000;
        mem[873] = 16'b0101101010000000;
        mem[874] = 16'b0101101011000000;
        mem[875] = 16'b0101101100000000;
        mem[876] = 16'b0101101101000000;
        mem[877] = 16'b0101101110000000;
        mem[878] = 16'b0101101111000000;
        mem[879] = 16'b0101110000000000;
        mem[880] = 16'b0101110001000000;
        mem[881] = 16'b0101110010000000;
        mem[882] = 16'b0101110011000000;
        mem[883] = 16'b0101110100000000;
        mem[884] = 16'b0101110101000000;
        mem[885] = 16'b0101110110000000;
        mem[886] = 16'b0101110111000000;
        mem[887] = 16'b0101111000000000;
        mem[888] = 16'b0101111001000000;
        mem[889] = 16'b0101111010000000;
        mem[890] = 16'b0101111011000000;
        mem[891] = 16'b0101111100000000;
        mem[892] = 16'b0101111101000000;
        mem[893] = 16'b0101111110000000;
        mem[894] = 16'b0101111111000000;
        mem[895] = 16'b0110000000000000;
        mem[896] = 16'b0110000001000000;
        mem[897] = 16'b0110000010000000;
        mem[898] = 16'b0110000011000000;
        mem[899] = 16'b0110000100000000;
        mem[900] = 16'b0110000101000000;
        mem[901] = 16'b0110000110000000;
        mem[902] = 16'b0110000111000000;
        mem[903] = 16'b0110001000000000;
        mem[904] = 16'b0110001001000000;
        mem[905] = 16'b0110001010000000;
        mem[906] = 16'b0110001011000000;
        mem[907] = 16'b0110001100000000;
        mem[908] = 16'b0110001101000000;
        mem[909] = 16'b0110001110000000;
        mem[910] = 16'b0110001111000000;
        mem[911] = 16'b0110010000000000;
        mem[912] = 16'b0110010001000000;
        mem[913] = 16'b0110010010000000;
        mem[914] = 16'b0110010011000000;
        mem[915] = 16'b0110010100000000;
        mem[916] = 16'b0110010101000000;
        mem[917] = 16'b0110010110000000;
        mem[918] = 16'b0110010111000000;
        mem[919] = 16'b0110011000000000;
        mem[920] = 16'b0110011001000000;
        mem[921] = 16'b0110011010000000;
        mem[922] = 16'b0110011011000000;
        mem[923] = 16'b0110011100000000;
        mem[924] = 16'b0110011101000000;
        mem[925] = 16'b0110011110000000;
        mem[926] = 16'b0110011111000000;
        mem[927] = 16'b0110100000000000;
        mem[928] = 16'b0110100001000000;
        mem[929] = 16'b0110100010000000;
        mem[930] = 16'b0110100011000000;
        mem[931] = 16'b0110100100000000;
        mem[932] = 16'b0110100101000000;
        mem[933] = 16'b0110100110000000;
        mem[934] = 16'b0110100111000000;
        mem[935] = 16'b0110101000000000;
        mem[936] = 16'b0110101001000000;
        mem[937] = 16'b0110101010000000;
        mem[938] = 16'b0110101011000000;
        mem[939] = 16'b0110101100000000;
        mem[940] = 16'b0110101101000000;
        mem[941] = 16'b0110101110000000;
        mem[942] = 16'b0110101111000000;
        mem[943] = 16'b0110110000000000;
        mem[944] = 16'b0110110001000000;
        mem[945] = 16'b0110110010000000;
        mem[946] = 16'b0110110011000000;
        mem[947] = 16'b0110110100000000;
        mem[948] = 16'b0110110101000000;
        mem[949] = 16'b0110110110000000;
        mem[950] = 16'b0110110111000000;
        mem[951] = 16'b0110111000000000;
        mem[952] = 16'b0110111001000000;
        mem[953] = 16'b0110111010000000;
        mem[954] = 16'b0110111011000000;
        mem[955] = 16'b0110111100000000;
        mem[956] = 16'b0110111101000000;
        mem[957] = 16'b0110111110000000;
        mem[958] = 16'b0110111111000000;
        mem[959] = 16'b0111000000000000;
        mem[960] = 16'b0111000001000000;
        mem[961] = 16'b0111000010000000;
        mem[962] = 16'b0111000011000000;
        mem[963] = 16'b0111000100000000;
        mem[964] = 16'b0111000101000000;
        mem[965] = 16'b0111000110000000;
        mem[966] = 16'b0111000111000000;
        mem[967] = 16'b0111001000000000;
        mem[968] = 16'b0111001001000000;
        mem[969] = 16'b0111001010000000;
        mem[970] = 16'b0111001011000000;
        mem[971] = 16'b0111001100000000;
        mem[972] = 16'b0111001101000000;
        mem[973] = 16'b0111001110000000;
        mem[974] = 16'b0111001111000000;
        mem[975] = 16'b0111010000000000;
        mem[976] = 16'b0111010001000000;
        mem[977] = 16'b0111010010000000;
        mem[978] = 16'b0111010011000000;
        mem[979] = 16'b0111010100000000;
        mem[980] = 16'b0111010101000000;
        mem[981] = 16'b0111010110000000;
        mem[982] = 16'b0111010111000000;
        mem[983] = 16'b0111011000000000;
        mem[984] = 16'b0111011001000000;
        mem[985] = 16'b0111011010000000;
        mem[986] = 16'b0111011011000000;
        mem[987] = 16'b0111011100000000;
        mem[988] = 16'b0111011101000000;
        mem[989] = 16'b0111011110000000;
        mem[990] = 16'b0111011111000000;
        mem[991] = 16'b0111100000000000;
        mem[992] = 16'b0111100001000000;
        mem[993] = 16'b0111100010000000;
        mem[994] = 16'b0111100011000000;
        mem[995] = 16'b0111100100000000;
        mem[996] = 16'b0111100101000000;
        mem[997] = 16'b0111100110000000;
        mem[998] = 16'b0111100111000000;
        mem[999] = 16'b0111101000000000;
        mem[1000] = 16'b0111101001000000;
        mem[1001] = 16'b0111101010000000;
        mem[1002] = 16'b0111101011000000;
        mem[1003] = 16'b0111101100000000;
        mem[1004] = 16'b0111101101000000;
        mem[1005] = 16'b0111101110000000;
        mem[1006] = 16'b0111101111000000;
        mem[1007] = 16'b0111110000000000;
        mem[1008] = 16'b0111110001000000;
        mem[1009] = 16'b0111110010000000;
        mem[1010] = 16'b0111110011000000;
        mem[1011] = 16'b0111110100000000;
        mem[1012] = 16'b0111110101000000;
        mem[1013] = 16'b0111110110000000;
        mem[1014] = 16'b0111110111000000;
        mem[1015] = 16'b0111111000000000;
        mem[1016] = 16'b0111111001000000;
        mem[1017] = 16'b0111111010000000;
        mem[1018] = 16'b0111111011000000;
        mem[1019] = 16'b0111111100000000;
        mem[1020] = 16'b0111111101000000;
        mem[1021] = 16'b0111111110000000;
        mem[1022] = 16'b0111111111000000;
    end
endmodule