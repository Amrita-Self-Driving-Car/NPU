//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.08.2021 22:17:08
// Design Name: 
// Module Name: X_Rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module X_Rom(
  input load_mem
);
    reg [31:0] mem [511:0];
    always @(posedge load_mem)
    begin
        mem[0] = 10'b1100000001;
        mem[1] = 10'b1100000010;
        mem[2] = 10'b1100000011;
        mem[3] = 10'b1100000100;
        mem[4] = 10'b1100000101;
        mem[5] = 10'b1100000110;
        mem[6] = 10'b1100000111;
        mem[7] = 10'b1100001000;
        mem[8] = 10'b1100001001;
        mem[9] = 10'b1100001010;
        mem[10] = 10'b1100001011;
        mem[11] = 10'b1100001100;
        mem[12] = 10'b1100001101;
        mem[13] = 10'b1100001110;
        mem[14] = 10'b1100001111;
        mem[15] = 10'b1100010000;
        mem[16] = 10'b1100010001;
        mem[17] = 10'b1100010010;
        mem[18] = 10'b1100010011;
        mem[19] = 10'b1100010100;
        mem[20] = 10'b1100010101;
        mem[21] = 10'b1100010110;
        mem[22] = 10'b1100010111;
        mem[23] = 10'b1100011000;
        mem[24] = 10'b1100011001;
        mem[25] = 10'b1100011010;
        mem[26] = 10'b1100011011;
        mem[27] = 10'b1100011100;
        mem[28] = 10'b1100011101;
        mem[29] = 10'b1100011110;
        mem[30] = 10'b1100011111;
        mem[31] = 10'b1100100000;
        mem[32] = 10'b1100100001;
        mem[33] = 10'b1100100010;
        mem[34] = 10'b1100100011;
        mem[35] = 10'b1100100100;
        mem[36] = 10'b1100100101;
        mem[37] = 10'b1100100110;
        mem[38] = 10'b1100100111;
        mem[39] = 10'b1100101000;
        mem[40] = 10'b1100101001;
        mem[41] = 10'b1100101010;
        mem[42] = 10'b1100101011;
        mem[43] = 10'b1100101100;
        mem[44] = 10'b1100101101;
        mem[45] = 10'b1100101110;
        mem[46] = 10'b1100101111;
        mem[47] = 10'b1100110000;
        mem[48] = 10'b1100110001;
        mem[49] = 10'b1100110010;
        mem[50] = 10'b1100110011;
        mem[51] = 10'b1100110100;
        mem[52] = 10'b1100110101;
        mem[53] = 10'b1100110110;
        mem[54] = 10'b1100110111;
        mem[55] = 10'b1100111000;
        mem[56] = 10'b1100111001;
        mem[57] = 10'b1100111010;
        mem[58] = 10'b1100111011;
        mem[59] = 10'b1100111100;
        mem[60] = 10'b1100111101;
        mem[61] = 10'b1100111110;
        mem[62] = 10'b1100111111;
        mem[63] = 10'b1101000000;
        mem[64] = 10'b1101000001;
        mem[65] = 10'b1101000010;
        mem[66] = 10'b1101000011;
        mem[67] = 10'b1101000100;
        mem[68] = 10'b1101000101;
        mem[69] = 10'b1101000110;
        mem[70] = 10'b1101000111;
        mem[71] = 10'b1101001000;
        mem[72] = 10'b1101001001;
        mem[73] = 10'b1101001010;
        mem[74] = 10'b1101001011;
        mem[75] = 10'b1101001100;
        mem[76] = 10'b1101001101;
        mem[77] = 10'b1101001110;
        mem[78] = 10'b1101001111;
        mem[79] = 10'b1101010000;
        mem[80] = 10'b1101010001;
        mem[81] = 10'b1101010010;
        mem[82] = 10'b1101010011;
        mem[83] = 10'b1101010100;
        mem[84] = 10'b1101010101;
        mem[85] = 10'b1101010110;
        mem[86] = 10'b1101010111;
        mem[87] = 10'b1101011000;
        mem[88] = 10'b1101011001;
        mem[89] = 10'b1101011010;
        mem[90] = 10'b1101011011;
        mem[91] = 10'b1101011100;
        mem[92] = 10'b1101011101;
        mem[93] = 10'b1101011110;
        mem[94] = 10'b1101011111;
        mem[95] = 10'b1101100000;
        mem[96] = 10'b1101100001;
        mem[97] = 10'b1101100010;
        mem[98] = 10'b1101100011;
        mem[99] = 10'b1101100100;
        mem[100] = 10'b1101100101;
        mem[101] = 10'b1101100110;
        mem[102] = 10'b1101100111;
        mem[103] = 10'b1101101000;
        mem[104] = 10'b1101101001;
        mem[105] = 10'b1101101010;
        mem[106] = 10'b1101101011;
        mem[107] = 10'b1101101100;
        mem[108] = 10'b1101101101;
        mem[109] = 10'b1101101110;
        mem[110] = 10'b1101101111;
        mem[111] = 10'b1101110000;
        mem[112] = 10'b1101110001;
        mem[113] = 10'b1101110010;
        mem[114] = 10'b1101110011;
        mem[115] = 10'b1101110100;
        mem[116] = 10'b1101110101;
        mem[117] = 10'b1101110110;
        mem[118] = 10'b1101110111;
        mem[119] = 10'b1101111000;
        mem[120] = 10'b1101111001;
        mem[121] = 10'b1101111010;
        mem[122] = 10'b1101111011;
        mem[123] = 10'b1101111100;
        mem[124] = 10'b1101111101;
        mem[125] = 10'b1101111110;
        mem[126] = 10'b1101111111;
        mem[127] = 10'b1110000000;
        mem[128] = 10'b1110000001;
        mem[129] = 10'b1110000010;
        mem[130] = 10'b1110000011;
        mem[131] = 10'b1110000100;
        mem[132] = 10'b1110000101;
        mem[133] = 10'b1110000110;
        mem[134] = 10'b1110000111;
        mem[135] = 10'b1110001000;
        mem[136] = 10'b1110001001;
        mem[137] = 10'b1110001010;
        mem[138] = 10'b1110001011;
        mem[139] = 10'b1110001100;
        mem[140] = 10'b1110001101;
        mem[141] = 10'b1110001110;
        mem[142] = 10'b1110001111;
        mem[143] = 10'b1110010000;
        mem[144] = 10'b1110010001;
        mem[145] = 10'b1110010010;
        mem[146] = 10'b1110010011;
        mem[147] = 10'b1110010100;
        mem[148] = 10'b1110010101;
        mem[149] = 10'b1110010110;
        mem[150] = 10'b1110010111;
        mem[151] = 10'b1110011000;
        mem[152] = 10'b1110011001;
        mem[153] = 10'b1110011010;
        mem[154] = 10'b1110011011;
        mem[155] = 10'b1110011100;
        mem[156] = 10'b1110011101;
        mem[157] = 10'b1110011110;
        mem[158] = 10'b1110011111;
        mem[159] = 10'b1110100000;
        mem[160] = 10'b1110100001;
        mem[161] = 10'b1110100010;
        mem[162] = 10'b1110100011;
        mem[163] = 10'b1110100100;
        mem[164] = 10'b1110100101;
        mem[165] = 10'b1110100110;
        mem[166] = 10'b1110100111;
        mem[167] = 10'b1110101000;
        mem[168] = 10'b1110101001;
        mem[169] = 10'b1110101010;
        mem[170] = 10'b1110101011;
        mem[171] = 10'b1110101100;
        mem[172] = 10'b1110101101;
        mem[173] = 10'b1110101110;
        mem[174] = 10'b1110101111;
        mem[175] = 10'b1110110000;
        mem[176] = 10'b1110110001;
        mem[177] = 10'b1110110010;
        mem[178] = 10'b1110110011;
        mem[179] = 10'b1110110100;
        mem[180] = 10'b1110110101;
        mem[181] = 10'b1110110110;
        mem[182] = 10'b1110110111;
        mem[183] = 10'b1110111000;
        mem[184] = 10'b1110111001;
        mem[185] = 10'b1110111010;
        mem[186] = 10'b1110111011;
        mem[187] = 10'b1110111100;
        mem[188] = 10'b1110111101;
        mem[189] = 10'b1110111110;
        mem[190] = 10'b1110111111;
        mem[191] = 10'b1111000000;
        mem[192] = 10'b1111000001;
        mem[193] = 10'b1111000010;
        mem[194] = 10'b1111000011;
        mem[195] = 10'b1111000100;
        mem[196] = 10'b1111000101;
        mem[197] = 10'b1111000110;
        mem[198] = 10'b1111000111;
        mem[199] = 10'b1111001000;
        mem[200] = 10'b1111001001;
        mem[201] = 10'b1111001010;
        mem[202] = 10'b1111001011;
        mem[203] = 10'b1111001100;
        mem[204] = 10'b1111001101;
        mem[205] = 10'b1111001110;
        mem[206] = 10'b1111001111;
        mem[207] = 10'b1111010000;
        mem[208] = 10'b1111010001;
        mem[209] = 10'b1111010010;
        mem[210] = 10'b1111010011;
        mem[211] = 10'b1111010100;
        mem[212] = 10'b1111010101;
        mem[213] = 10'b1111010110;
        mem[214] = 10'b1111010111;
        mem[215] = 10'b1111011000;
        mem[216] = 10'b1111011001;
        mem[217] = 10'b1111011010;
        mem[218] = 10'b1111011011;
        mem[219] = 10'b1111011100;
        mem[220] = 10'b1111011101;
        mem[221] = 10'b1111011110;
        mem[222] = 10'b1111011111;
        mem[223] = 10'b1111100000;
        mem[224] = 10'b1111100001;
        mem[225] = 10'b1111100010;
        mem[226] = 10'b1111100011;
        mem[227] = 10'b1111100100;
        mem[228] = 10'b1111100101;
        mem[229] = 10'b1111100110;
        mem[230] = 10'b1111100111;
        mem[231] = 10'b1111101000;
        mem[232] = 10'b1111101001;
        mem[233] = 10'b1111101010;
        mem[234] = 10'b1111101011;
        mem[235] = 10'b1111101100;
        mem[236] = 10'b1111101101;
        mem[237] = 10'b1111101110;
        mem[238] = 10'b1111101111;
        mem[239] = 10'b1111110000;
        mem[240] = 10'b1111110001;
        mem[241] = 10'b1111110010;
        mem[242] = 10'b1111110011;
        mem[243] = 10'b1111110100;
        mem[244] = 10'b1111110101;
        mem[245] = 10'b1111110110;
        mem[246] = 10'b1111110111;
        mem[247] = 10'b1111111000;
        mem[248] = 10'b1111111001;
        mem[249] = 10'b1111111010;
        mem[250] = 10'b1111111011;
        mem[251] = 10'b1111111100;
        mem[252] = 10'b1111111101;
        mem[253] = 10'b1111111110;
        mem[254] = 10'b1111111111;
        mem[255] = 10'b0000000000;
        mem[256] = 10'b0000000001;
        mem[257] = 10'b0000000010;
        mem[258] = 10'b0000000011;
        mem[259] = 10'b0000000100;
        mem[260] = 10'b0000000101;
        mem[261] = 10'b0000000110;
        mem[262] = 10'b0000000111;
        mem[263] = 10'b0000001000;
        mem[264] = 10'b0000001001;
        mem[265] = 10'b0000001010;
        mem[266] = 10'b0000001011;
        mem[267] = 10'b0000001100;
        mem[268] = 10'b0000001101;
        mem[269] = 10'b0000001110;
        mem[270] = 10'b0000001111;
        mem[271] = 10'b0000010000;
        mem[272] = 10'b0000010001;
        mem[273] = 10'b0000010010;
        mem[274] = 10'b0000010011;
        mem[275] = 10'b0000010100;
        mem[276] = 10'b0000010101;
        mem[277] = 10'b0000010110;
        mem[278] = 10'b0000010111;
        mem[279] = 10'b0000011000;
        mem[280] = 10'b0000011001;
        mem[281] = 10'b0000011010;
        mem[282] = 10'b0000011011;
        mem[283] = 10'b0000011100;
        mem[284] = 10'b0000011101;
        mem[285] = 10'b0000011110;
        mem[286] = 10'b0000011111;
        mem[287] = 10'b0000100000;
        mem[288] = 10'b0000100001;
        mem[289] = 10'b0000100010;
        mem[290] = 10'b0000100011;
        mem[291] = 10'b0000100100;
        mem[292] = 10'b0000100101;
        mem[293] = 10'b0000100110;
        mem[294] = 10'b0000100111;
        mem[295] = 10'b0000101000;
        mem[296] = 10'b0000101001;
        mem[297] = 10'b0000101010;
        mem[298] = 10'b0000101011;
        mem[299] = 10'b0000101100;
        mem[300] = 10'b0000101101;
        mem[301] = 10'b0000101110;
        mem[302] = 10'b0000101111;
        mem[303] = 10'b0000110000;
        mem[304] = 10'b0000110001;
        mem[305] = 10'b0000110010;
        mem[306] = 10'b0000110011;
        mem[307] = 10'b0000110100;
        mem[308] = 10'b0000110101;
        mem[309] = 10'b0000110110;
        mem[310] = 10'b0000110111;
        mem[311] = 10'b0000111000;
        mem[312] = 10'b0000111001;
        mem[313] = 10'b0000111010;
        mem[314] = 10'b0000111011;
        mem[315] = 10'b0000111100;
        mem[316] = 10'b0000111101;
        mem[317] = 10'b0000111110;
        mem[318] = 10'b0000111111;
        mem[319] = 10'b0001000000;
        mem[320] = 10'b0001000001;
        mem[321] = 10'b0001000010;
        mem[322] = 10'b0001000011;
        mem[323] = 10'b0001000100;
        mem[324] = 10'b0001000101;
        mem[325] = 10'b0001000110;
        mem[326] = 10'b0001000111;
        mem[327] = 10'b0001001000;
        mem[328] = 10'b0001001001;
        mem[329] = 10'b0001001010;
        mem[330] = 10'b0001001011;
        mem[331] = 10'b0001001100;
        mem[332] = 10'b0001001101;
        mem[333] = 10'b0001001110;
        mem[334] = 10'b0001001111;
        mem[335] = 10'b0001010000;
        mem[336] = 10'b0001010001;
        mem[337] = 10'b0001010010;
        mem[338] = 10'b0001010011;
        mem[339] = 10'b0001010100;
        mem[340] = 10'b0001010101;
        mem[341] = 10'b0001010110;
        mem[342] = 10'b0001010111;
        mem[343] = 10'b0001011000;
        mem[344] = 10'b0001011001;
        mem[345] = 10'b0001011010;
        mem[346] = 10'b0001011011;
        mem[347] = 10'b0001011100;
        mem[348] = 10'b0001011101;
        mem[349] = 10'b0001011110;
        mem[350] = 10'b0001011111;
        mem[351] = 10'b0001100000;
        mem[352] = 10'b0001100001;
        mem[353] = 10'b0001100010;
        mem[354] = 10'b0001100011;
        mem[355] = 10'b0001100100;
        mem[356] = 10'b0001100101;
        mem[357] = 10'b0001100110;
        mem[358] = 10'b0001100111;
        mem[359] = 10'b0001101000;
        mem[360] = 10'b0001101001;
        mem[361] = 10'b0001101010;
        mem[362] = 10'b0001101011;
        mem[363] = 10'b0001101100;
        mem[364] = 10'b0001101101;
        mem[365] = 10'b0001101110;
        mem[366] = 10'b0001101111;
        mem[367] = 10'b0001110000;
        mem[368] = 10'b0001110001;
        mem[369] = 10'b0001110010;
        mem[370] = 10'b0001110011;
        mem[371] = 10'b0001110100;
        mem[372] = 10'b0001110101;
        mem[373] = 10'b0001110110;
        mem[374] = 10'b0001110111;
        mem[375] = 10'b0001111000;
        mem[376] = 10'b0001111001;
        mem[377] = 10'b0001111010;
        mem[378] = 10'b0001111011;
        mem[379] = 10'b0001111100;
        mem[380] = 10'b0001111101;
        mem[381] = 10'b0001111110;
        mem[382] = 10'b0001111111;
        mem[383] = 10'b0010000000;
        mem[384] = 10'b0010000001;
        mem[385] = 10'b0010000010;
        mem[386] = 10'b0010000011;
        mem[387] = 10'b0010000100;
        mem[388] = 10'b0010000101;
        mem[389] = 10'b0010000110;
        mem[390] = 10'b0010000111;
        mem[391] = 10'b0010001000;
        mem[392] = 10'b0010001001;
        mem[393] = 10'b0010001010;
        mem[394] = 10'b0010001011;
        mem[395] = 10'b0010001100;
        mem[396] = 10'b0010001101;
        mem[397] = 10'b0010001110;
        mem[398] = 10'b0010001111;
        mem[399] = 10'b0010010000;
        mem[400] = 10'b0010010001;
        mem[401] = 10'b0010010010;
        mem[402] = 10'b0010010011;
        mem[403] = 10'b0010010100;
        mem[404] = 10'b0010010101;
        mem[405] = 10'b0010010110;
        mem[406] = 10'b0010010111;
        mem[407] = 10'b0010011000;
        mem[408] = 10'b0010011001;
        mem[409] = 10'b0010011010;
        mem[410] = 10'b0010011011;
        mem[411] = 10'b0010011100;
        mem[412] = 10'b0010011101;
        mem[413] = 10'b0010011110;
        mem[414] = 10'b0010011111;
        mem[415] = 10'b0010100000;
        mem[416] = 10'b0010100001;
        mem[417] = 10'b0010100010;
        mem[418] = 10'b0010100011;
        mem[419] = 10'b0010100100;
        mem[420] = 10'b0010100101;
        mem[421] = 10'b0010100110;
        mem[422] = 10'b0010100111;
        mem[423] = 10'b0010101000;
        mem[424] = 10'b0010101001;
        mem[425] = 10'b0010101010;
        mem[426] = 10'b0010101011;
        mem[427] = 10'b0010101100;
        mem[428] = 10'b0010101101;
        mem[429] = 10'b0010101110;
        mem[430] = 10'b0010101111;
        mem[431] = 10'b0010110000;
        mem[432] = 10'b0010110001;
        mem[433] = 10'b0010110010;
        mem[434] = 10'b0010110011;
        mem[435] = 10'b0010110100;
        mem[436] = 10'b0010110101;
        mem[437] = 10'b0010110110;
        mem[438] = 10'b0010110111;
        mem[439] = 10'b0010111000;
        mem[440] = 10'b0010111001;
        mem[441] = 10'b0010111010;
        mem[442] = 10'b0010111011;
        mem[443] = 10'b0010111100;
        mem[444] = 10'b0010111101;
        mem[445] = 10'b0010111110;
        mem[446] = 10'b0010111111;
        mem[447] = 10'b0011000000;
        mem[448] = 10'b0011000001;
        mem[449] = 10'b0011000010;
        mem[450] = 10'b0011000011;
        mem[451] = 10'b0011000100;
        mem[452] = 10'b0011000101;
        mem[453] = 10'b0011000110;
        mem[454] = 10'b0011000111;
        mem[455] = 10'b0011001000;
        mem[456] = 10'b0011001001;
        mem[457] = 10'b0011001010;
        mem[458] = 10'b0011001011;
        mem[459] = 10'b0011001100;
        mem[460] = 10'b0011001101;
        mem[461] = 10'b0011001110;
        mem[462] = 10'b0011001111;
        mem[463] = 10'b0011010000;
        mem[464] = 10'b0011010001;
        mem[465] = 10'b0011010010;
        mem[466] = 10'b0011010011;
        mem[467] = 10'b0011010100;
        mem[468] = 10'b0011010101;
        mem[469] = 10'b0011010110;
        mem[470] = 10'b0011010111;
        mem[471] = 10'b0011011000;
        mem[472] = 10'b0011011001;
        mem[473] = 10'b0011011010;
        mem[474] = 10'b0011011011;
        mem[475] = 10'b0011011100;
        mem[476] = 10'b0011011101;
        mem[477] = 10'b0011011110;
        mem[478] = 10'b0011011111;
        mem[479] = 10'b0011100000;
        mem[480] = 10'b0011100001;
        mem[481] = 10'b0011100010;
        mem[482] = 10'b0011100011;
        mem[483] = 10'b0011100100;
        mem[484] = 10'b0011100101;
        mem[485] = 10'b0011100110;
        mem[486] = 10'b0011100111;
        mem[487] = 10'b0011101000;
        mem[488] = 10'b0011101001;
        mem[489] = 10'b0011101010;
        mem[490] = 10'b0011101011;
        mem[491] = 10'b0011101100;
        mem[492] = 10'b0011101101;
        mem[493] = 10'b0011101110;
        mem[494] = 10'b0011101111;
        mem[495] = 10'b0011110000;
        mem[496] = 10'b0011110001;
        mem[497] = 10'b0011110010;
        mem[498] = 10'b0011110011;
        mem[499] = 10'b0011110100;
        mem[500] = 10'b0011110101;
        mem[501] = 10'b0011110110;
        mem[502] = 10'b0011110111;
        mem[503] = 10'b0011111000;
        mem[504] = 10'b0011111001;
        mem[505] = 10'b0011111010;
        mem[506] = 10'b0011111011;
        mem[507] = 10'b0011111100;
        mem[508] = 10'b0011111101;
        mem[509] = 10'b0011111110;
        mem[510] = 10'b0011111111;
    end
endmodule